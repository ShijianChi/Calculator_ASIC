
module mux4_1_0 ( selector, data_in_00, data_in_01, data_in_10, data_in_11, 
        data_out );
  input [1:0] selector;
  input [31:0] data_in_00;
  input [31:0] data_in_01;
  input [31:0] data_in_10;
  input [31:0] data_in_11;
  output [31:0] data_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  NOR2X2TS U1 ( .A(selector[0]), .B(selector[1]), .Y(n25) );
  NOR2BX1TS U2 ( .AN(selector[1]), .B(selector[0]), .Y(n29) );
  CLKBUFX2TS U3 ( .A(n29), .Y(n23) );
  NOR2BX1TS U4 ( .AN(selector[0]), .B(selector[1]), .Y(n26) );
  CLKBUFX2TS U5 ( .A(n26), .Y(n27) );
  AOI222XLTS U6 ( .A0(n23), .A1(data_in_10[6]), .B0(n27), .B1(data_in_01[6]), 
        .C0(n25), .C1(data_in_00[6]), .Y(n1) );
  INVX2TS U7 ( .A(n1), .Y(data_out[6]) );
  AOI222XLTS U8 ( .A0(n23), .A1(data_in_10[9]), .B0(n27), .B1(data_in_01[9]), 
        .C0(n25), .C1(data_in_00[9]), .Y(n2) );
  INVX2TS U9 ( .A(n2), .Y(data_out[9]) );
  AOI222XLTS U10 ( .A0(n23), .A1(data_in_10[1]), .B0(n27), .B1(data_in_01[1]), 
        .C0(n25), .C1(data_in_00[1]), .Y(n3) );
  INVX2TS U11 ( .A(n3), .Y(data_out[1]) );
  AOI222XLTS U12 ( .A0(n23), .A1(data_in_10[10]), .B0(n27), .B1(data_in_01[10]), .C0(n25), .C1(data_in_00[10]), .Y(n4) );
  INVX2TS U13 ( .A(n4), .Y(data_out[10]) );
  AOI222XLTS U14 ( .A0(n23), .A1(data_in_10[12]), .B0(n27), .B1(data_in_01[12]), .C0(n25), .C1(data_in_00[12]), .Y(n5) );
  INVX2TS U15 ( .A(n5), .Y(data_out[12]) );
  AOI222XLTS U16 ( .A0(n23), .A1(data_in_10[2]), .B0(n27), .B1(data_in_01[2]), 
        .C0(n25), .C1(data_in_00[2]), .Y(n6) );
  INVX2TS U17 ( .A(n6), .Y(data_out[2]) );
  AOI222XLTS U18 ( .A0(n23), .A1(data_in_10[16]), .B0(n27), .B1(data_in_01[16]), .C0(n25), .C1(data_in_00[16]), .Y(n7) );
  INVX2TS U19 ( .A(n7), .Y(data_out[16]) );
  AOI222XLTS U20 ( .A0(n23), .A1(data_in_10[4]), .B0(n27), .B1(data_in_01[4]), 
        .C0(n25), .C1(data_in_00[4]), .Y(n8) );
  INVX2TS U21 ( .A(n8), .Y(data_out[4]) );
  AOI222XLTS U22 ( .A0(n23), .A1(data_in_10[13]), .B0(n27), .B1(data_in_01[13]), .C0(n25), .C1(data_in_00[13]), .Y(n9) );
  INVX2TS U23 ( .A(n9), .Y(data_out[13]) );
  AOI222XLTS U24 ( .A0(n23), .A1(data_in_10[14]), .B0(n27), .B1(data_in_01[14]), .C0(n25), .C1(data_in_00[14]), .Y(n10) );
  INVX2TS U25 ( .A(n10), .Y(data_out[14]) );
  AOI222XLTS U26 ( .A0(n23), .A1(data_in_10[11]), .B0(n27), .B1(data_in_01[11]), .C0(n25), .C1(data_in_00[11]), .Y(n11) );
  INVX2TS U27 ( .A(n11), .Y(data_out[11]) );
  AOI222XLTS U28 ( .A0(n23), .A1(data_in_10[5]), .B0(n27), .B1(data_in_01[5]), 
        .C0(n25), .C1(data_in_00[5]), .Y(n12) );
  INVX2TS U29 ( .A(n12), .Y(data_out[5]) );
  AOI222XLTS U30 ( .A0(n23), .A1(data_in_10[3]), .B0(n27), .B1(data_in_01[3]), 
        .C0(n25), .C1(data_in_00[3]), .Y(n13) );
  INVX2TS U31 ( .A(n13), .Y(data_out[3]) );
  AOI222XLTS U32 ( .A0(n23), .A1(data_in_10[15]), .B0(n27), .B1(data_in_01[15]), .C0(n25), .C1(data_in_00[15]), .Y(n14) );
  INVX2TS U33 ( .A(n14), .Y(data_out[15]) );
  AOI222XLTS U34 ( .A0(n23), .A1(data_in_10[7]), .B0(n27), .B1(data_in_01[7]), 
        .C0(n25), .C1(data_in_00[7]), .Y(n15) );
  INVX2TS U35 ( .A(n15), .Y(data_out[7]) );
  AOI222XLTS U36 ( .A0(n23), .A1(data_in_10[8]), .B0(n27), .B1(data_in_01[8]), 
        .C0(n25), .C1(data_in_00[8]), .Y(n16) );
  INVX2TS U37 ( .A(n16), .Y(data_out[8]) );
  AOI222XLTS U38 ( .A0(n23), .A1(data_in_10[20]), .B0(n27), .B1(data_in_01[20]), .C0(n25), .C1(data_in_00[20]), .Y(n17) );
  INVX2TS U39 ( .A(n17), .Y(data_out[20]) );
  AOI222XLTS U40 ( .A0(n23), .A1(data_in_10[21]), .B0(n27), .B1(data_in_01[21]), .C0(n25), .C1(data_in_00[21]), .Y(n18) );
  INVX2TS U41 ( .A(n18), .Y(data_out[21]) );
  AOI222XLTS U42 ( .A0(n23), .A1(data_in_10[0]), .B0(n27), .B1(data_in_01[0]), 
        .C0(n25), .C1(data_in_00[0]), .Y(n19) );
  INVX2TS U43 ( .A(n19), .Y(data_out[0]) );
  AOI222XLTS U44 ( .A0(n23), .A1(data_in_10[22]), .B0(n27), .B1(data_in_01[22]), .C0(n25), .C1(data_in_00[22]), .Y(n20) );
  INVX2TS U45 ( .A(n20), .Y(data_out[22]) );
  AOI222XLTS U46 ( .A0(n23), .A1(data_in_10[18]), .B0(n27), .B1(data_in_01[18]), .C0(n25), .C1(data_in_00[18]), .Y(n21) );
  INVX2TS U47 ( .A(n21), .Y(data_out[18]) );
  AOI222XLTS U48 ( .A0(n23), .A1(data_in_10[19]), .B0(n27), .B1(data_in_01[19]), .C0(n25), .C1(data_in_00[19]), .Y(n22) );
  INVX2TS U49 ( .A(n22), .Y(data_out[19]) );
  AOI222XLTS U50 ( .A0(n23), .A1(data_in_10[17]), .B0(n27), .B1(data_in_01[17]), .C0(n25), .C1(data_in_00[17]), .Y(n24) );
  INVX2TS U51 ( .A(n24), .Y(data_out[17]) );
  AO22XLTS U52 ( .A0(n27), .A1(data_in_01[24]), .B0(n25), .B1(data_in_00[24]), 
        .Y(data_out[24]) );
  AO22XLTS U53 ( .A0(n27), .A1(data_in_01[25]), .B0(n25), .B1(data_in_00[25]), 
        .Y(data_out[25]) );
  AO22XLTS U54 ( .A0(n27), .A1(data_in_01[26]), .B0(n25), .B1(data_in_00[26]), 
        .Y(data_out[26]) );
  AO22XLTS U55 ( .A0(n27), .A1(data_in_01[27]), .B0(n25), .B1(data_in_00[27]), 
        .Y(data_out[27]) );
  AO22XLTS U56 ( .A0(n27), .A1(data_in_01[28]), .B0(n25), .B1(data_in_00[28]), 
        .Y(data_out[28]) );
  AO22XLTS U57 ( .A0(n26), .A1(data_in_01[29]), .B0(n25), .B1(data_in_00[29]), 
        .Y(data_out[29]) );
  AO22XLTS U58 ( .A0(n26), .A1(data_in_01[30]), .B0(n25), .B1(data_in_00[30]), 
        .Y(data_out[30]) );
  AO22XLTS U59 ( .A0(n26), .A1(data_in_01[31]), .B0(n25), .B1(data_in_00[31]), 
        .Y(data_out[31]) );
  AOI22X1TS U60 ( .A0(n27), .A1(data_in_01[23]), .B0(n25), .B1(data_in_00[23]), 
        .Y(n28) );
  NAND2BXLTS U61 ( .AN(n29), .B(n28), .Y(data_out[23]) );
endmodule


module mux2_1_0 ( selector, data_in_0, data_in_1, data_out );
  input [31:0] data_in_0;
  input [31:0] data_in_1;
  output [31:0] data_out;
  input selector;
  wire   n1;

  INVX2TS U1 ( .A(selector), .Y(n1) );
  NAND2BXLTS U2 ( .AN(data_in_0[23]), .B(n1), .Y(data_out[23]) );
  CLKAND2X2TS U3 ( .A(data_in_0[24]), .B(n1), .Y(data_out[24]) );
  CLKAND2X2TS U4 ( .A(data_in_0[25]), .B(n1), .Y(data_out[25]) );
  CLKAND2X2TS U5 ( .A(data_in_0[26]), .B(n1), .Y(data_out[26]) );
  CLKAND2X2TS U6 ( .A(data_in_0[27]), .B(n1), .Y(data_out[27]) );
  CLKAND2X2TS U7 ( .A(data_in_0[28]), .B(n1), .Y(data_out[28]) );
  CLKAND2X2TS U8 ( .A(data_in_0[29]), .B(n1), .Y(data_out[29]) );
  CLKAND2X2TS U9 ( .A(data_in_0[30]), .B(n1), .Y(data_out[30]) );
  CLKAND2X2TS U10 ( .A(data_in_0[31]), .B(n1), .Y(data_out[31]) );
  AO22XLTS U11 ( .A0(selector), .A1(data_in_1[0]), .B0(n1), .B1(data_in_0[0]), 
        .Y(data_out[0]) );
  AO22XLTS U12 ( .A0(selector), .A1(data_in_1[1]), .B0(n1), .B1(data_in_0[1]), 
        .Y(data_out[1]) );
  AO22XLTS U13 ( .A0(selector), .A1(data_in_1[2]), .B0(n1), .B1(data_in_0[2]), 
        .Y(data_out[2]) );
  AO22XLTS U14 ( .A0(selector), .A1(data_in_1[3]), .B0(n1), .B1(data_in_0[3]), 
        .Y(data_out[3]) );
  AO22XLTS U15 ( .A0(selector), .A1(data_in_1[4]), .B0(n1), .B1(data_in_0[4]), 
        .Y(data_out[4]) );
  AO22XLTS U16 ( .A0(selector), .A1(data_in_1[5]), .B0(n1), .B1(data_in_0[5]), 
        .Y(data_out[5]) );
  AO22XLTS U17 ( .A0(selector), .A1(data_in_1[6]), .B0(n1), .B1(data_in_0[6]), 
        .Y(data_out[6]) );
  AO22XLTS U18 ( .A0(selector), .A1(data_in_1[7]), .B0(n1), .B1(data_in_0[7]), 
        .Y(data_out[7]) );
  AO22XLTS U19 ( .A0(selector), .A1(data_in_1[8]), .B0(n1), .B1(data_in_0[8]), 
        .Y(data_out[8]) );
  AO22XLTS U20 ( .A0(selector), .A1(data_in_1[9]), .B0(n1), .B1(data_in_0[9]), 
        .Y(data_out[9]) );
  AO22XLTS U21 ( .A0(selector), .A1(data_in_1[10]), .B0(n1), .B1(data_in_0[10]), .Y(data_out[10]) );
  AO22XLTS U22 ( .A0(selector), .A1(data_in_1[11]), .B0(n1), .B1(data_in_0[11]), .Y(data_out[11]) );
  AO22XLTS U23 ( .A0(selector), .A1(data_in_1[12]), .B0(n1), .B1(data_in_0[12]), .Y(data_out[12]) );
  AO22XLTS U24 ( .A0(selector), .A1(data_in_1[13]), .B0(n1), .B1(data_in_0[13]), .Y(data_out[13]) );
  AO22XLTS U25 ( .A0(selector), .A1(data_in_1[14]), .B0(n1), .B1(data_in_0[14]), .Y(data_out[14]) );
  AO22XLTS U26 ( .A0(selector), .A1(data_in_1[15]), .B0(n1), .B1(data_in_0[15]), .Y(data_out[15]) );
  AO22XLTS U27 ( .A0(selector), .A1(data_in_1[16]), .B0(n1), .B1(data_in_0[16]), .Y(data_out[16]) );
  AO22XLTS U28 ( .A0(selector), .A1(data_in_1[17]), .B0(n1), .B1(data_in_0[17]), .Y(data_out[17]) );
  AO22XLTS U29 ( .A0(selector), .A1(data_in_1[18]), .B0(n1), .B1(data_in_0[18]), .Y(data_out[18]) );
  AO22XLTS U30 ( .A0(selector), .A1(data_in_1[19]), .B0(n1), .B1(data_in_0[19]), .Y(data_out[19]) );
  AO22XLTS U31 ( .A0(selector), .A1(data_in_1[20]), .B0(n1), .B1(data_in_0[20]), .Y(data_out[20]) );
  AO22XLTS U32 ( .A0(selector), .A1(data_in_1[21]), .B0(n1), .B1(data_in_0[21]), .Y(data_out[21]) );
  AO22XLTS U33 ( .A0(selector), .A1(data_in_1[22]), .B0(n1), .B1(data_in_0[22]), .Y(data_out[22]) );
endmodule


module register_0 ( clk, load, data_in, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, load;


  EDFFX1TS \data_out_buffer_reg[31]  ( .D(data_in[31]), .E(load), .CK(clk), 
        .Q(data_out[31]) );
  EDFFX1TS \data_out_buffer_reg[30]  ( .D(data_in[30]), .E(load), .CK(clk), 
        .Q(data_out[30]) );
  EDFFX1TS \data_out_buffer_reg[29]  ( .D(data_in[29]), .E(load), .CK(clk), 
        .Q(data_out[29]) );
  EDFFX1TS \data_out_buffer_reg[28]  ( .D(data_in[28]), .E(load), .CK(clk), 
        .Q(data_out[28]) );
  EDFFX1TS \data_out_buffer_reg[27]  ( .D(data_in[27]), .E(load), .CK(clk), 
        .Q(data_out[27]) );
  EDFFX1TS \data_out_buffer_reg[26]  ( .D(data_in[26]), .E(load), .CK(clk), 
        .Q(data_out[26]) );
  EDFFX1TS \data_out_buffer_reg[25]  ( .D(data_in[25]), .E(load), .CK(clk), 
        .Q(data_out[25]) );
  EDFFX1TS \data_out_buffer_reg[24]  ( .D(data_in[24]), .E(load), .CK(clk), 
        .Q(data_out[24]) );
  EDFFX1TS \data_out_buffer_reg[23]  ( .D(data_in[23]), .E(load), .CK(clk), 
        .Q(data_out[23]) );
  EDFFX1TS \data_out_buffer_reg[22]  ( .D(data_in[22]), .E(load), .CK(clk), 
        .Q(data_out[22]) );
  EDFFX1TS \data_out_buffer_reg[21]  ( .D(data_in[21]), .E(load), .CK(clk), 
        .Q(data_out[21]) );
  EDFFX1TS \data_out_buffer_reg[20]  ( .D(data_in[20]), .E(load), .CK(clk), 
        .Q(data_out[20]) );
  EDFFX1TS \data_out_buffer_reg[19]  ( .D(data_in[19]), .E(load), .CK(clk), 
        .Q(data_out[19]) );
  EDFFX1TS \data_out_buffer_reg[18]  ( .D(data_in[18]), .E(load), .CK(clk), 
        .Q(data_out[18]) );
  EDFFX1TS \data_out_buffer_reg[17]  ( .D(data_in[17]), .E(load), .CK(clk), 
        .Q(data_out[17]) );
  EDFFX1TS \data_out_buffer_reg[16]  ( .D(data_in[16]), .E(load), .CK(clk), 
        .Q(data_out[16]) );
  EDFFX1TS \data_out_buffer_reg[15]  ( .D(data_in[15]), .E(load), .CK(clk), 
        .Q(data_out[15]) );
  EDFFX1TS \data_out_buffer_reg[14]  ( .D(data_in[14]), .E(load), .CK(clk), 
        .Q(data_out[14]) );
  EDFFX1TS \data_out_buffer_reg[13]  ( .D(data_in[13]), .E(load), .CK(clk), 
        .Q(data_out[13]) );
  EDFFX1TS \data_out_buffer_reg[12]  ( .D(data_in[12]), .E(load), .CK(clk), 
        .Q(data_out[12]) );
  EDFFX1TS \data_out_buffer_reg[11]  ( .D(data_in[11]), .E(load), .CK(clk), 
        .Q(data_out[11]) );
  EDFFX1TS \data_out_buffer_reg[10]  ( .D(data_in[10]), .E(load), .CK(clk), 
        .Q(data_out[10]) );
  EDFFX1TS \data_out_buffer_reg[9]  ( .D(data_in[9]), .E(load), .CK(clk), .Q(
        data_out[9]) );
  EDFFX1TS \data_out_buffer_reg[8]  ( .D(data_in[8]), .E(load), .CK(clk), .Q(
        data_out[8]) );
  EDFFX1TS \data_out_buffer_reg[7]  ( .D(data_in[7]), .E(load), .CK(clk), .Q(
        data_out[7]) );
  EDFFX1TS \data_out_buffer_reg[6]  ( .D(data_in[6]), .E(load), .CK(clk), .Q(
        data_out[6]) );
  EDFFX1TS \data_out_buffer_reg[5]  ( .D(data_in[5]), .E(load), .CK(clk), .Q(
        data_out[5]) );
  EDFFX1TS \data_out_buffer_reg[4]  ( .D(data_in[4]), .E(load), .CK(clk), .Q(
        data_out[4]) );
  EDFFX1TS \data_out_buffer_reg[3]  ( .D(data_in[3]), .E(load), .CK(clk), .Q(
        data_out[3]) );
  EDFFX1TS \data_out_buffer_reg[2]  ( .D(data_in[2]), .E(load), .CK(clk), .Q(
        data_out[2]) );
  EDFFX1TS \data_out_buffer_reg[1]  ( .D(data_in[1]), .E(load), .CK(clk), .Q(
        data_out[1]) );
  EDFFX1TS \data_out_buffer_reg[0]  ( .D(data_in[0]), .E(load), .CK(clk), .Q(
        data_out[0]) );
endmodule


module mult32_0 ( A, B, Product );
  input [31:0] A;
  input [31:0] B;
  output [63:0] Product;
  wire   \mult_x_1/n1250 , \mult_x_1/n1249 , \mult_x_1/n1248 ,
         \mult_x_1/n1247 , \mult_x_1/n1246 , \mult_x_1/n1245 ,
         \mult_x_1/n1244 , \mult_x_1/n1243 , \mult_x_1/n1242 ,
         \mult_x_1/n1241 , \mult_x_1/n1240 , \mult_x_1/n1239 ,
         \mult_x_1/n1238 , \mult_x_1/n1237 , \mult_x_1/n1236 ,
         \mult_x_1/n1235 , \mult_x_1/n1234 , \mult_x_1/n1233 ,
         \mult_x_1/n1232 , \mult_x_1/n1231 , \mult_x_1/n1230 ,
         \mult_x_1/n1229 , \mult_x_1/n1228 , \mult_x_1/n1227 ,
         \mult_x_1/n1226 , \mult_x_1/n1225 , \mult_x_1/n1224 ,
         \mult_x_1/n1223 , \mult_x_1/n1218 , \mult_x_1/n1217 ,
         \mult_x_1/n1216 , \mult_x_1/n1215 , \mult_x_1/n1214 ,
         \mult_x_1/n1213 , \mult_x_1/n1212 , \mult_x_1/n1211 ,
         \mult_x_1/n1210 , \mult_x_1/n1209 , \mult_x_1/n1208 ,
         \mult_x_1/n1207 , \mult_x_1/n1206 , \mult_x_1/n1205 ,
         \mult_x_1/n1204 , \mult_x_1/n1203 , \mult_x_1/n1202 ,
         \mult_x_1/n1201 , \mult_x_1/n1200 , \mult_x_1/n1199 ,
         \mult_x_1/n1198 , \mult_x_1/n1197 , \mult_x_1/n1196 ,
         \mult_x_1/n1195 , \mult_x_1/n1194 , \mult_x_1/n1193 ,
         \mult_x_1/n1192 , \mult_x_1/n1191 , \mult_x_1/n1190 ,
         \mult_x_1/n1189 , \mult_x_1/n1188 , \mult_x_1/n1180 ,
         \mult_x_1/n1179 , \mult_x_1/n1178 , \mult_x_1/n1177 ,
         \mult_x_1/n1176 , \mult_x_1/n1175 , \mult_x_1/n1174 ,
         \mult_x_1/n1173 , \mult_x_1/n1172 , \mult_x_1/n1171 ,
         \mult_x_1/n1170 , \mult_x_1/n1169 , \mult_x_1/n1168 ,
         \mult_x_1/n1167 , \mult_x_1/n1166 , \mult_x_1/n1165 ,
         \mult_x_1/n1164 , \mult_x_1/n1163 , \mult_x_1/n1162 ,
         \mult_x_1/n1161 , \mult_x_1/n1160 , \mult_x_1/n1159 ,
         \mult_x_1/n1158 , \mult_x_1/n1157 , \mult_x_1/n1156 ,
         \mult_x_1/n1155 , \mult_x_1/n1154 , \mult_x_1/n1153 ,
         \mult_x_1/n1148 , \mult_x_1/n1147 , \mult_x_1/n1146 ,
         \mult_x_1/n1145 , \mult_x_1/n1144 , \mult_x_1/n1143 ,
         \mult_x_1/n1142 , \mult_x_1/n1141 , \mult_x_1/n1140 ,
         \mult_x_1/n1139 , \mult_x_1/n1138 , \mult_x_1/n1137 ,
         \mult_x_1/n1136 , \mult_x_1/n1135 , \mult_x_1/n1134 ,
         \mult_x_1/n1133 , \mult_x_1/n1132 , \mult_x_1/n1131 ,
         \mult_x_1/n1130 , \mult_x_1/n1129 , \mult_x_1/n1128 ,
         \mult_x_1/n1127 , \mult_x_1/n1126 , \mult_x_1/n1125 ,
         \mult_x_1/n1124 , \mult_x_1/n1123 , \mult_x_1/n1122 ,
         \mult_x_1/n1121 , \mult_x_1/n1120 , \mult_x_1/n1119 ,
         \mult_x_1/n1118 , \mult_x_1/n1110 , \mult_x_1/n1109 ,
         \mult_x_1/n1108 , \mult_x_1/n1107 , \mult_x_1/n1106 ,
         \mult_x_1/n1105 , \mult_x_1/n1104 , \mult_x_1/n1103 ,
         \mult_x_1/n1102 , \mult_x_1/n1101 , \mult_x_1/n1100 ,
         \mult_x_1/n1099 , \mult_x_1/n1098 , \mult_x_1/n1097 ,
         \mult_x_1/n1096 , \mult_x_1/n1095 , \mult_x_1/n1094 ,
         \mult_x_1/n1093 , \mult_x_1/n1092 , \mult_x_1/n1091 ,
         \mult_x_1/n1090 , \mult_x_1/n1089 , \mult_x_1/n1088 ,
         \mult_x_1/n1087 , \mult_x_1/n1086 , \mult_x_1/n1085 ,
         \mult_x_1/n1084 , \mult_x_1/n1083 , \mult_x_1/n1078 ,
         \mult_x_1/n1077 , \mult_x_1/n1076 , \mult_x_1/n1075 ,
         \mult_x_1/n1074 , \mult_x_1/n1073 , \mult_x_1/n1072 ,
         \mult_x_1/n1071 , \mult_x_1/n1070 , \mult_x_1/n1069 ,
         \mult_x_1/n1068 , \mult_x_1/n1067 , \mult_x_1/n1066 ,
         \mult_x_1/n1065 , \mult_x_1/n1064 , \mult_x_1/n1063 ,
         \mult_x_1/n1062 , \mult_x_1/n1061 , \mult_x_1/n1060 ,
         \mult_x_1/n1059 , \mult_x_1/n1058 , \mult_x_1/n1057 ,
         \mult_x_1/n1056 , \mult_x_1/n1055 , \mult_x_1/n1054 ,
         \mult_x_1/n1053 , \mult_x_1/n1052 , \mult_x_1/n1051 ,
         \mult_x_1/n1050 , \mult_x_1/n1049 , \mult_x_1/n1048 ,
         \mult_x_1/n1040 , \mult_x_1/n1039 , \mult_x_1/n1038 ,
         \mult_x_1/n1037 , \mult_x_1/n1036 , \mult_x_1/n1035 ,
         \mult_x_1/n1034 , \mult_x_1/n1033 , \mult_x_1/n1032 ,
         \mult_x_1/n1031 , \mult_x_1/n1030 , \mult_x_1/n1029 ,
         \mult_x_1/n1028 , \mult_x_1/n1027 , \mult_x_1/n1026 ,
         \mult_x_1/n1025 , \mult_x_1/n1024 , \mult_x_1/n1023 ,
         \mult_x_1/n1022 , \mult_x_1/n1021 , \mult_x_1/n1020 ,
         \mult_x_1/n1019 , \mult_x_1/n1018 , \mult_x_1/n1017 ,
         \mult_x_1/n1016 , \mult_x_1/n1015 , \mult_x_1/n1014 ,
         \mult_x_1/n1013 , \mult_x_1/n1008 , \mult_x_1/n1007 ,
         \mult_x_1/n1006 , \mult_x_1/n1005 , \mult_x_1/n1004 ,
         \mult_x_1/n1003 , \mult_x_1/n1002 , \mult_x_1/n1001 ,
         \mult_x_1/n1000 , \mult_x_1/n999 , \mult_x_1/n998 , \mult_x_1/n997 ,
         \mult_x_1/n996 , \mult_x_1/n995 , \mult_x_1/n994 , \mult_x_1/n993 ,
         \mult_x_1/n992 , \mult_x_1/n991 , \mult_x_1/n990 , \mult_x_1/n989 ,
         \mult_x_1/n988 , \mult_x_1/n987 , \mult_x_1/n986 , \mult_x_1/n985 ,
         \mult_x_1/n984 , \mult_x_1/n983 , \mult_x_1/n982 , \mult_x_1/n981 ,
         \mult_x_1/n980 , \mult_x_1/n979 , \mult_x_1/n978 , \mult_x_1/n966 ,
         \mult_x_1/n965 , \mult_x_1/n964 , \mult_x_1/n963 , \mult_x_1/n960 ,
         \mult_x_1/n959 , \mult_x_1/n958 , \mult_x_1/n957 , \mult_x_1/n954 ,
         \mult_x_1/n953 , \mult_x_1/n952 , \mult_x_1/n951 , \mult_x_1/n949 ,
         \mult_x_1/n948 , \mult_x_1/n947 , \mult_x_1/n946 , \mult_x_1/n945 ,
         \mult_x_1/n933 , \mult_x_1/n932 , \mult_x_1/n928 , \mult_x_1/n927 ,
         \mult_x_1/n923 , \mult_x_1/n922 , \mult_x_1/n918 , \mult_x_1/n917 ,
         \mult_x_1/n916 , \mult_x_1/n798 , \mult_x_1/n796 , \mult_x_1/n795 ,
         \mult_x_1/n793 , \mult_x_1/n792 , \mult_x_1/n791 , \mult_x_1/n790 ,
         \mult_x_1/n788 , \mult_x_1/n787 , \mult_x_1/n786 , \mult_x_1/n785 ,
         \mult_x_1/n783 , \mult_x_1/n782 , \mult_x_1/n781 , \mult_x_1/n778 ,
         \mult_x_1/n776 , \mult_x_1/n775 , \mult_x_1/n774 , \mult_x_1/n771 ,
         \mult_x_1/n769 , \mult_x_1/n768 , \mult_x_1/n767 , \mult_x_1/n765 ,
         \mult_x_1/n764 , \mult_x_1/n763 , \mult_x_1/n762 , \mult_x_1/n761 ,
         \mult_x_1/n760 , \mult_x_1/n759 , \mult_x_1/n757 , \mult_x_1/n756 ,
         \mult_x_1/n755 , \mult_x_1/n754 , \mult_x_1/n753 , \mult_x_1/n752 ,
         \mult_x_1/n751 , \mult_x_1/n749 , \mult_x_1/n748 , \mult_x_1/n747 ,
         \mult_x_1/n746 , \mult_x_1/n745 , \mult_x_1/n744 , \mult_x_1/n743 ,
         \mult_x_1/n741 , \mult_x_1/n740 , \mult_x_1/n739 , \mult_x_1/n738 ,
         \mult_x_1/n737 , \mult_x_1/n736 , \mult_x_1/n733 , \mult_x_1/n731 ,
         \mult_x_1/n730 , \mult_x_1/n729 , \mult_x_1/n728 , \mult_x_1/n727 ,
         \mult_x_1/n726 , \mult_x_1/n723 , \mult_x_1/n721 , \mult_x_1/n720 ,
         \mult_x_1/n719 , \mult_x_1/n718 , \mult_x_1/n717 , \mult_x_1/n716 ,
         \mult_x_1/n714 , \mult_x_1/n713 , \mult_x_1/n712 , \mult_x_1/n711 ,
         \mult_x_1/n710 , \mult_x_1/n709 , \mult_x_1/n708 , \mult_x_1/n707 ,
         \mult_x_1/n706 , \mult_x_1/n705 , \mult_x_1/n703 , \mult_x_1/n702 ,
         \mult_x_1/n701 , \mult_x_1/n700 , \mult_x_1/n699 , \mult_x_1/n698 ,
         \mult_x_1/n697 , \mult_x_1/n696 , \mult_x_1/n695 , \mult_x_1/n694 ,
         \mult_x_1/n692 , \mult_x_1/n691 , \mult_x_1/n690 , \mult_x_1/n689 ,
         \mult_x_1/n688 , \mult_x_1/n687 , \mult_x_1/n686 , \mult_x_1/n685 ,
         \mult_x_1/n684 , \mult_x_1/n683 , \mult_x_1/n681 , \mult_x_1/n680 ,
         \mult_x_1/n679 , \mult_x_1/n678 , \mult_x_1/n677 , \mult_x_1/n676 ,
         \mult_x_1/n675 , \mult_x_1/n674 , \mult_x_1/n673 , \mult_x_1/n670 ,
         \mult_x_1/n668 , \mult_x_1/n667 , \mult_x_1/n666 , \mult_x_1/n665 ,
         \mult_x_1/n664 , \mult_x_1/n663 , \mult_x_1/n662 , \mult_x_1/n661 ,
         \mult_x_1/n660 , \mult_x_1/n657 , \mult_x_1/n655 , \mult_x_1/n654 ,
         \mult_x_1/n653 , \mult_x_1/n652 , \mult_x_1/n651 , \mult_x_1/n650 ,
         \mult_x_1/n649 , \mult_x_1/n648 , \mult_x_1/n647 , \mult_x_1/n645 ,
         \mult_x_1/n644 , \mult_x_1/n643 , \mult_x_1/n642 , \mult_x_1/n641 ,
         \mult_x_1/n640 , \mult_x_1/n639 , \mult_x_1/n638 , \mult_x_1/n637 ,
         \mult_x_1/n636 , \mult_x_1/n635 , \mult_x_1/n634 , \mult_x_1/n633 ,
         \mult_x_1/n631 , \mult_x_1/n630 , \mult_x_1/n629 , \mult_x_1/n628 ,
         \mult_x_1/n627 , \mult_x_1/n626 , \mult_x_1/n625 , \mult_x_1/n624 ,
         \mult_x_1/n623 , \mult_x_1/n622 , \mult_x_1/n621 , \mult_x_1/n620 ,
         \mult_x_1/n619 , \mult_x_1/n617 , \mult_x_1/n616 , \mult_x_1/n615 ,
         \mult_x_1/n614 , \mult_x_1/n613 , \mult_x_1/n612 , \mult_x_1/n611 ,
         \mult_x_1/n610 , \mult_x_1/n609 , \mult_x_1/n608 , \mult_x_1/n607 ,
         \mult_x_1/n606 , \mult_x_1/n605 , \mult_x_1/n603 , \mult_x_1/n602 ,
         \mult_x_1/n601 , \mult_x_1/n600 , \mult_x_1/n599 , \mult_x_1/n598 ,
         \mult_x_1/n597 , \mult_x_1/n596 , \mult_x_1/n595 , \mult_x_1/n594 ,
         \mult_x_1/n593 , \mult_x_1/n592 , \mult_x_1/n591 , \mult_x_1/n589 ,
         \mult_x_1/n588 , \mult_x_1/n587 , \mult_x_1/n586 , \mult_x_1/n585 ,
         \mult_x_1/n584 , \mult_x_1/n583 , \mult_x_1/n582 , \mult_x_1/n581 ,
         \mult_x_1/n580 , \mult_x_1/n579 , \mult_x_1/n578 , \mult_x_1/n577 ,
         \mult_x_1/n575 , \mult_x_1/n574 , \mult_x_1/n573 , \mult_x_1/n572 ,
         \mult_x_1/n571 , \mult_x_1/n570 , \mult_x_1/n569 , \mult_x_1/n568 ,
         \mult_x_1/n567 , \mult_x_1/n566 , \mult_x_1/n565 , \mult_x_1/n564 ,
         \mult_x_1/n563 , \mult_x_1/n561 , \mult_x_1/n560 , \mult_x_1/n559 ,
         \mult_x_1/n558 , \mult_x_1/n557 , \mult_x_1/n556 , \mult_x_1/n555 ,
         \mult_x_1/n554 , \mult_x_1/n553 , \mult_x_1/n552 , \mult_x_1/n551 ,
         \mult_x_1/n550 , \mult_x_1/n549 , \mult_x_1/n548 , \mult_x_1/n547 ,
         \mult_x_1/n546 , \mult_x_1/n545 , \mult_x_1/n544 , \mult_x_1/n543 ,
         \mult_x_1/n542 , \mult_x_1/n541 , \mult_x_1/n540 , \mult_x_1/n539 ,
         \mult_x_1/n538 , \mult_x_1/n537 , \mult_x_1/n536 , \mult_x_1/n535 ,
         \mult_x_1/n534 , \mult_x_1/n533 , \mult_x_1/n532 , \mult_x_1/n531 ,
         \mult_x_1/n530 , \mult_x_1/n529 , \mult_x_1/n528 , \mult_x_1/n527 ,
         \mult_x_1/n526 , \mult_x_1/n525 , \mult_x_1/n524 , \mult_x_1/n523 ,
         \mult_x_1/n522 , \mult_x_1/n521 , \mult_x_1/n520 , \mult_x_1/n519 ,
         \mult_x_1/n518 , \mult_x_1/n517 , \mult_x_1/n516 , \mult_x_1/n515 ,
         \mult_x_1/n514 , \mult_x_1/n513 , \mult_x_1/n512 , \mult_x_1/n511 ,
         \mult_x_1/n510 , \mult_x_1/n509 , \mult_x_1/n508 , \mult_x_1/n507 ,
         \mult_x_1/n506 , \mult_x_1/n505 , \mult_x_1/n504 , \mult_x_1/n503 ,
         \mult_x_1/n502 , \mult_x_1/n501 , \mult_x_1/n500 , \mult_x_1/n499 ,
         \mult_x_1/n498 , \mult_x_1/n497 , \mult_x_1/n496 , \mult_x_1/n495 ,
         \mult_x_1/n494 , \mult_x_1/n493 , \mult_x_1/n492 , \mult_x_1/n491 ,
         \mult_x_1/n490 , \mult_x_1/n489 , \mult_x_1/n488 , \mult_x_1/n487 ,
         \mult_x_1/n486 , \mult_x_1/n485 , \mult_x_1/n484 , \mult_x_1/n483 ,
         \mult_x_1/n482 , \mult_x_1/n481 , \mult_x_1/n480 , \mult_x_1/n479 ,
         \mult_x_1/n478 , \mult_x_1/n477 , \mult_x_1/n476 , \mult_x_1/n475 ,
         \mult_x_1/n474 , \mult_x_1/n473 , \mult_x_1/n472 , \mult_x_1/n471 ,
         \mult_x_1/n470 , \mult_x_1/n469 , \mult_x_1/n468 , \mult_x_1/n467 ,
         \mult_x_1/n465 , \mult_x_1/n464 , \mult_x_1/n463 , \mult_x_1/n462 ,
         \mult_x_1/n461 , \mult_x_1/n460 , \mult_x_1/n459 , \mult_x_1/n458 ,
         \mult_x_1/n457 , \mult_x_1/n456 , \mult_x_1/n455 , \mult_x_1/n454 ,
         \mult_x_1/n453 , \mult_x_1/n452 , \mult_x_1/n451 , \mult_x_1/n450 ,
         \mult_x_1/n449 , \mult_x_1/n448 , \mult_x_1/n447 , \mult_x_1/n446 ,
         \mult_x_1/n445 , \mult_x_1/n444 , \mult_x_1/n443 , \mult_x_1/n442 ,
         \mult_x_1/n440 , \mult_x_1/n439 , \mult_x_1/n438 , \mult_x_1/n437 ,
         \mult_x_1/n436 , \mult_x_1/n435 , \mult_x_1/n434 , \mult_x_1/n433 ,
         \mult_x_1/n432 , \mult_x_1/n431 , \mult_x_1/n430 , \mult_x_1/n428 ,
         \mult_x_1/n427 , \mult_x_1/n426 , \mult_x_1/n425 , \mult_x_1/n424 ,
         \mult_x_1/n423 , \mult_x_1/n422 , \mult_x_1/n421 , \mult_x_1/n420 ,
         \mult_x_1/n419 , \mult_x_1/n418 , \mult_x_1/n417 , \mult_x_1/n416 ,
         \mult_x_1/n415 , \mult_x_1/n414 , \mult_x_1/n413 , \mult_x_1/n412 ,
         \mult_x_1/n411 , \mult_x_1/n410 , \mult_x_1/n409 , \mult_x_1/n408 ,
         \mult_x_1/n407 , \mult_x_1/n406 , \mult_x_1/n405 , \mult_x_1/n404 ,
         \mult_x_1/n403 , \mult_x_1/n402 , \mult_x_1/n401 , \mult_x_1/n400 ,
         \mult_x_1/n399 , \mult_x_1/n398 , \mult_x_1/n397 , \mult_x_1/n396 ,
         \mult_x_1/n394 , \mult_x_1/n393 , \mult_x_1/n392 , \mult_x_1/n391 ,
         \mult_x_1/n390 , \mult_x_1/n389 , \mult_x_1/n388 , \mult_x_1/n387 ,
         \mult_x_1/n386 , \mult_x_1/n385 , \mult_x_1/n384 , \mult_x_1/n383 ,
         \mult_x_1/n382 , \mult_x_1/n381 , \mult_x_1/n380 , \mult_x_1/n379 ,
         \mult_x_1/n378 , \mult_x_1/n377 , \mult_x_1/n375 , \mult_x_1/n374 ,
         \mult_x_1/n373 , \mult_x_1/n372 , \mult_x_1/n371 , \mult_x_1/n370 ,
         \mult_x_1/n369 , \mult_x_1/n368 , \mult_x_1/n366 , \mult_x_1/n365 ,
         \mult_x_1/n364 , \mult_x_1/n363 , \mult_x_1/n362 , \mult_x_1/n361 ,
         \mult_x_1/n360 , \mult_x_1/n359 , \mult_x_1/n358 , \mult_x_1/n357 ,
         \mult_x_1/n356 , \mult_x_1/n355 , \mult_x_1/n354 , \mult_x_1/n353 ,
         \mult_x_1/n352 , \mult_x_1/n351 , \mult_x_1/n350 , \mult_x_1/n349 ,
         \mult_x_1/n348 , \mult_x_1/n347 , \mult_x_1/n346 , \mult_x_1/n345 ,
         \mult_x_1/n344 , \mult_x_1/n343 , \mult_x_1/n341 , \mult_x_1/n340 ,
         \mult_x_1/n339 , \mult_x_1/n338 , \mult_x_1/n337 , \mult_x_1/n336 ,
         \mult_x_1/n335 , \mult_x_1/n334 , \mult_x_1/n333 , \mult_x_1/n332 ,
         \mult_x_1/n331 , \mult_x_1/n330 , \mult_x_1/n328 , \mult_x_1/n326 ,
         \mult_x_1/n325 , \mult_x_1/n324 , \mult_x_1/n322 , \mult_x_1/n321 ,
         \mult_x_1/n320 , \mult_x_1/n319 , \mult_x_1/n318 , \mult_x_1/n317 ,
         \mult_x_1/n316 , \mult_x_1/n315 , \mult_x_1/n314 , \mult_x_1/n313 ,
         \mult_x_1/n312 , \mult_x_1/n311 , \mult_x_1/n310 , \mult_x_1/n309 ,
         \mult_x_1/n307 , \mult_x_1/n306 , \mult_x_1/n305 , \mult_x_1/n304 ,
         \mult_x_1/n303 , \mult_x_1/n302 , \mult_x_1/n297 , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674;

  CMPR42X1TS \mult_x_1/U485  ( .A(\mult_x_1/n795 ), .B(\mult_x_1/n1218 ), .C(
        \mult_x_1/n798 ), .D(\mult_x_1/n1250 ), .ICI(\mult_x_1/n796 ), .S(
        \mult_x_1/n793 ), .ICO(\mult_x_1/n791 ), .CO(\mult_x_1/n792 ) );
  CMPR42X1TS \mult_x_1/U483  ( .A(\mult_x_1/n790 ), .B(\mult_x_1/n1217 ), .C(
        \mult_x_1/n791 ), .D(\mult_x_1/n1249 ), .ICI(\mult_x_1/n792 ), .S(
        \mult_x_1/n788 ), .ICO(\mult_x_1/n786 ), .CO(\mult_x_1/n787 ) );
  CMPR42X1TS \mult_x_1/U481  ( .A(\mult_x_1/n785 ), .B(\mult_x_1/n1216 ), .C(
        \mult_x_1/n786 ), .D(\mult_x_1/n1248 ), .ICI(\mult_x_1/n787 ), .S(
        \mult_x_1/n783 ), .ICO(\mult_x_1/n781 ), .CO(\mult_x_1/n782 ) );
  CMPR42X1TS \mult_x_1/U478  ( .A(\mult_x_1/n778 ), .B(\mult_x_1/n781 ), .C(
        \mult_x_1/n1215 ), .D(\mult_x_1/n1247 ), .ICI(\mult_x_1/n782 ), .S(
        \mult_x_1/n776 ), .ICO(\mult_x_1/n774 ), .CO(\mult_x_1/n775 ) );
  CMPR42X1TS \mult_x_1/U475  ( .A(\mult_x_1/n771 ), .B(\mult_x_1/n774 ), .C(
        \mult_x_1/n1214 ), .D(\mult_x_1/n1246 ), .ICI(\mult_x_1/n775 ), .S(
        \mult_x_1/n769 ), .ICO(\mult_x_1/n767 ), .CO(\mult_x_1/n768 ) );
  CMPR42X1TS \mult_x_1/U472  ( .A(\mult_x_1/n764 ), .B(\mult_x_1/n767 ), .C(
        \mult_x_1/n1213 ), .D(\mult_x_1/n1245 ), .ICI(\mult_x_1/n768 ), .S(
        \mult_x_1/n762 ), .ICO(\mult_x_1/n760 ), .CO(\mult_x_1/n761 ) );
  CMPR42X1TS \mult_x_1/U470  ( .A(\mult_x_1/n759 ), .B(\mult_x_1/n1148 ), .C(
        \mult_x_1/n765 ), .D(\mult_x_1/n1180 ), .ICI(\mult_x_1/n763 ), .S(
        \mult_x_1/n757 ), .ICO(\mult_x_1/n755 ), .CO(\mult_x_1/n756 ) );
  CMPR42X1TS \mult_x_1/U469  ( .A(\mult_x_1/n757 ), .B(\mult_x_1/n760 ), .C(
        \mult_x_1/n1212 ), .D(\mult_x_1/n1244 ), .ICI(\mult_x_1/n761 ), .S(
        \mult_x_1/n754 ), .ICO(\mult_x_1/n752 ), .CO(\mult_x_1/n753 ) );
  CMPR42X1TS \mult_x_1/U467  ( .A(\mult_x_1/n751 ), .B(\mult_x_1/n1147 ), .C(
        \mult_x_1/n755 ), .D(\mult_x_1/n1179 ), .ICI(\mult_x_1/n756 ), .S(
        \mult_x_1/n749 ), .ICO(\mult_x_1/n747 ), .CO(\mult_x_1/n748 ) );
  CMPR42X1TS \mult_x_1/U466  ( .A(\mult_x_1/n749 ), .B(\mult_x_1/n752 ), .C(
        \mult_x_1/n1211 ), .D(\mult_x_1/n1243 ), .ICI(\mult_x_1/n753 ), .S(
        \mult_x_1/n746 ), .ICO(\mult_x_1/n744 ), .CO(\mult_x_1/n745 ) );
  CMPR42X1TS \mult_x_1/U464  ( .A(\mult_x_1/n743 ), .B(\mult_x_1/n1146 ), .C(
        \mult_x_1/n747 ), .D(\mult_x_1/n1178 ), .ICI(\mult_x_1/n748 ), .S(
        \mult_x_1/n741 ), .ICO(\mult_x_1/n739 ), .CO(\mult_x_1/n740 ) );
  CMPR42X1TS \mult_x_1/U463  ( .A(\mult_x_1/n741 ), .B(\mult_x_1/n744 ), .C(
        \mult_x_1/n1210 ), .D(\mult_x_1/n1242 ), .ICI(\mult_x_1/n745 ), .S(
        \mult_x_1/n738 ), .ICO(\mult_x_1/n736 ), .CO(\mult_x_1/n737 ) );
  CMPR42X1TS \mult_x_1/U460  ( .A(\mult_x_1/n733 ), .B(\mult_x_1/n739 ), .C(
        \mult_x_1/n1145 ), .D(\mult_x_1/n1177 ), .ICI(\mult_x_1/n740 ), .S(
        \mult_x_1/n731 ), .ICO(\mult_x_1/n729 ), .CO(\mult_x_1/n730 ) );
  CMPR42X1TS \mult_x_1/U459  ( .A(\mult_x_1/n731 ), .B(\mult_x_1/n736 ), .C(
        \mult_x_1/n1209 ), .D(\mult_x_1/n1241 ), .ICI(\mult_x_1/n737 ), .S(
        \mult_x_1/n728 ), .ICO(\mult_x_1/n726 ), .CO(\mult_x_1/n727 ) );
  CMPR42X1TS \mult_x_1/U456  ( .A(\mult_x_1/n723 ), .B(\mult_x_1/n729 ), .C(
        \mult_x_1/n1144 ), .D(\mult_x_1/n1176 ), .ICI(\mult_x_1/n730 ), .S(
        \mult_x_1/n721 ), .ICO(\mult_x_1/n719 ), .CO(\mult_x_1/n720 ) );
  CMPR42X1TS \mult_x_1/U455  ( .A(\mult_x_1/n721 ), .B(\mult_x_1/n726 ), .C(
        \mult_x_1/n1208 ), .D(\mult_x_1/n1240 ), .ICI(\mult_x_1/n727 ), .S(
        \mult_x_1/n718 ), .ICO(\mult_x_1/n716 ), .CO(\mult_x_1/n717 ) );
  CMPR42X1TS \mult_x_1/U452  ( .A(\mult_x_1/n713 ), .B(\mult_x_1/n719 ), .C(
        \mult_x_1/n1143 ), .D(\mult_x_1/n1175 ), .ICI(\mult_x_1/n720 ), .S(
        \mult_x_1/n711 ), .ICO(\mult_x_1/n709 ), .CO(\mult_x_1/n710 ) );
  CMPR42X1TS \mult_x_1/U451  ( .A(\mult_x_1/n711 ), .B(\mult_x_1/n716 ), .C(
        \mult_x_1/n1207 ), .D(\mult_x_1/n1239 ), .ICI(\mult_x_1/n717 ), .S(
        \mult_x_1/n708 ), .ICO(\mult_x_1/n706 ), .CO(\mult_x_1/n707 ) );
  CMPR42X1TS \mult_x_1/U449  ( .A(\mult_x_1/n705 ), .B(\mult_x_1/n1078 ), .C(
        \mult_x_1/n714 ), .D(\mult_x_1/n1110 ), .ICI(\mult_x_1/n712 ), .S(
        \mult_x_1/n703 ), .ICO(\mult_x_1/n701 ), .CO(\mult_x_1/n702 ) );
  CMPR42X1TS \mult_x_1/U448  ( .A(\mult_x_1/n703 ), .B(\mult_x_1/n709 ), .C(
        \mult_x_1/n1142 ), .D(\mult_x_1/n1174 ), .ICI(\mult_x_1/n710 ), .S(
        \mult_x_1/n700 ), .ICO(\mult_x_1/n698 ), .CO(\mult_x_1/n699 ) );
  CMPR42X1TS \mult_x_1/U447  ( .A(\mult_x_1/n700 ), .B(\mult_x_1/n706 ), .C(
        \mult_x_1/n1206 ), .D(\mult_x_1/n1238 ), .ICI(\mult_x_1/n707 ), .S(
        \mult_x_1/n697 ), .ICO(\mult_x_1/n695 ), .CO(\mult_x_1/n696 ) );
  CMPR42X1TS \mult_x_1/U445  ( .A(\mult_x_1/n694 ), .B(\mult_x_1/n1077 ), .C(
        \mult_x_1/n701 ), .D(\mult_x_1/n1109 ), .ICI(\mult_x_1/n702 ), .S(
        \mult_x_1/n692 ), .ICO(\mult_x_1/n690 ), .CO(\mult_x_1/n691 ) );
  CMPR42X1TS \mult_x_1/U444  ( .A(\mult_x_1/n692 ), .B(\mult_x_1/n698 ), .C(
        \mult_x_1/n1141 ), .D(\mult_x_1/n1173 ), .ICI(\mult_x_1/n699 ), .S(
        \mult_x_1/n689 ), .ICO(\mult_x_1/n687 ), .CO(\mult_x_1/n688 ) );
  CMPR42X1TS \mult_x_1/U443  ( .A(\mult_x_1/n689 ), .B(\mult_x_1/n695 ), .C(
        \mult_x_1/n1205 ), .D(\mult_x_1/n1237 ), .ICI(\mult_x_1/n696 ), .S(
        \mult_x_1/n686 ), .ICO(\mult_x_1/n684 ), .CO(\mult_x_1/n685 ) );
  CMPR42X1TS \mult_x_1/U441  ( .A(\mult_x_1/n683 ), .B(\mult_x_1/n1076 ), .C(
        \mult_x_1/n690 ), .D(\mult_x_1/n1108 ), .ICI(\mult_x_1/n691 ), .S(
        \mult_x_1/n681 ), .ICO(\mult_x_1/n679 ), .CO(\mult_x_1/n680 ) );
  CMPR42X1TS \mult_x_1/U440  ( .A(\mult_x_1/n681 ), .B(\mult_x_1/n687 ), .C(
        \mult_x_1/n1140 ), .D(\mult_x_1/n1172 ), .ICI(\mult_x_1/n688 ), .S(
        \mult_x_1/n678 ), .ICO(\mult_x_1/n676 ), .CO(\mult_x_1/n677 ) );
  CMPR42X1TS \mult_x_1/U439  ( .A(\mult_x_1/n678 ), .B(\mult_x_1/n684 ), .C(
        \mult_x_1/n1204 ), .D(\mult_x_1/n1236 ), .ICI(\mult_x_1/n685 ), .S(
        \mult_x_1/n675 ), .ICO(\mult_x_1/n673 ), .CO(\mult_x_1/n674 ) );
  CMPR42X1TS \mult_x_1/U436  ( .A(\mult_x_1/n670 ), .B(\mult_x_1/n679 ), .C(
        \mult_x_1/n1075 ), .D(\mult_x_1/n1107 ), .ICI(\mult_x_1/n680 ), .S(
        \mult_x_1/n668 ), .ICO(\mult_x_1/n666 ), .CO(\mult_x_1/n667 ) );
  CMPR42X1TS \mult_x_1/U435  ( .A(\mult_x_1/n668 ), .B(\mult_x_1/n676 ), .C(
        \mult_x_1/n1139 ), .D(\mult_x_1/n1171 ), .ICI(\mult_x_1/n677 ), .S(
        \mult_x_1/n665 ), .ICO(\mult_x_1/n663 ), .CO(\mult_x_1/n664 ) );
  CMPR42X1TS \mult_x_1/U434  ( .A(\mult_x_1/n665 ), .B(\mult_x_1/n673 ), .C(
        \mult_x_1/n1203 ), .D(\mult_x_1/n1235 ), .ICI(\mult_x_1/n674 ), .S(
        \mult_x_1/n662 ), .ICO(\mult_x_1/n660 ), .CO(\mult_x_1/n661 ) );
  CMPR42X1TS \mult_x_1/U431  ( .A(\mult_x_1/n657 ), .B(\mult_x_1/n666 ), .C(
        \mult_x_1/n1074 ), .D(\mult_x_1/n1106 ), .ICI(\mult_x_1/n667 ), .S(
        \mult_x_1/n655 ), .ICO(\mult_x_1/n653 ), .CO(\mult_x_1/n654 ) );
  CMPR42X1TS \mult_x_1/U430  ( .A(\mult_x_1/n655 ), .B(\mult_x_1/n663 ), .C(
        \mult_x_1/n1138 ), .D(\mult_x_1/n1170 ), .ICI(\mult_x_1/n664 ), .S(
        \mult_x_1/n652 ), .ICO(\mult_x_1/n650 ), .CO(\mult_x_1/n651 ) );
  CMPR42X1TS \mult_x_1/U429  ( .A(\mult_x_1/n652 ), .B(\mult_x_1/n660 ), .C(
        \mult_x_1/n1202 ), .D(\mult_x_1/n1234 ), .ICI(\mult_x_1/n661 ), .S(
        \mult_x_1/n649 ), .ICO(\mult_x_1/n647 ), .CO(\mult_x_1/n648 ) );
  CMPR42X1TS \mult_x_1/U426  ( .A(\mult_x_1/n644 ), .B(\mult_x_1/n653 ), .C(
        \mult_x_1/n1073 ), .D(\mult_x_1/n1105 ), .ICI(\mult_x_1/n654 ), .S(
        \mult_x_1/n642 ), .ICO(\mult_x_1/n640 ), .CO(\mult_x_1/n641 ) );
  CMPR42X1TS \mult_x_1/U425  ( .A(\mult_x_1/n642 ), .B(\mult_x_1/n650 ), .C(
        \mult_x_1/n1137 ), .D(\mult_x_1/n1169 ), .ICI(\mult_x_1/n651 ), .S(
        \mult_x_1/n639 ), .ICO(\mult_x_1/n637 ), .CO(\mult_x_1/n638 ) );
  CMPR42X1TS \mult_x_1/U424  ( .A(\mult_x_1/n639 ), .B(\mult_x_1/n647 ), .C(
        \mult_x_1/n1201 ), .D(\mult_x_1/n1233 ), .ICI(\mult_x_1/n648 ), .S(
        \mult_x_1/n636 ), .ICO(\mult_x_1/n634 ), .CO(\mult_x_1/n635 ) );
  CMPR42X1TS \mult_x_1/U422  ( .A(\mult_x_1/n633 ), .B(\mult_x_1/n1008 ), .C(
        \mult_x_1/n645 ), .D(\mult_x_1/n1040 ), .ICI(\mult_x_1/n643 ), .S(
        \mult_x_1/n631 ), .ICO(\mult_x_1/n629 ), .CO(\mult_x_1/n630 ) );
  CMPR42X1TS \mult_x_1/U421  ( .A(\mult_x_1/n631 ), .B(\mult_x_1/n640 ), .C(
        \mult_x_1/n1072 ), .D(\mult_x_1/n1104 ), .ICI(\mult_x_1/n641 ), .S(
        \mult_x_1/n628 ), .ICO(\mult_x_1/n626 ), .CO(\mult_x_1/n627 ) );
  CMPR42X1TS \mult_x_1/U420  ( .A(\mult_x_1/n628 ), .B(\mult_x_1/n637 ), .C(
        \mult_x_1/n1136 ), .D(\mult_x_1/n1168 ), .ICI(\mult_x_1/n638 ), .S(
        \mult_x_1/n625 ), .ICO(\mult_x_1/n623 ), .CO(\mult_x_1/n624 ) );
  CMPR42X1TS \mult_x_1/U419  ( .A(\mult_x_1/n625 ), .B(\mult_x_1/n634 ), .C(
        \mult_x_1/n1200 ), .D(\mult_x_1/n1232 ), .ICI(\mult_x_1/n635 ), .S(
        \mult_x_1/n622 ), .ICO(\mult_x_1/n620 ), .CO(\mult_x_1/n621 ) );
  CMPR42X1TS \mult_x_1/U417  ( .A(\mult_x_1/n619 ), .B(\mult_x_1/n1007 ), .C(
        \mult_x_1/n629 ), .D(\mult_x_1/n1039 ), .ICI(\mult_x_1/n630 ), .S(
        \mult_x_1/n617 ), .ICO(\mult_x_1/n615 ), .CO(\mult_x_1/n616 ) );
  CMPR42X1TS \mult_x_1/U416  ( .A(\mult_x_1/n617 ), .B(\mult_x_1/n626 ), .C(
        \mult_x_1/n1071 ), .D(\mult_x_1/n1103 ), .ICI(\mult_x_1/n627 ), .S(
        \mult_x_1/n614 ), .ICO(\mult_x_1/n612 ), .CO(\mult_x_1/n613 ) );
  CMPR42X1TS \mult_x_1/U415  ( .A(\mult_x_1/n614 ), .B(\mult_x_1/n623 ), .C(
        \mult_x_1/n1135 ), .D(\mult_x_1/n1167 ), .ICI(\mult_x_1/n624 ), .S(
        \mult_x_1/n611 ), .ICO(\mult_x_1/n609 ), .CO(\mult_x_1/n610 ) );
  CMPR42X1TS \mult_x_1/U414  ( .A(\mult_x_1/n611 ), .B(\mult_x_1/n620 ), .C(
        \mult_x_1/n1199 ), .D(\mult_x_1/n1231 ), .ICI(\mult_x_1/n621 ), .S(
        \mult_x_1/n608 ), .ICO(\mult_x_1/n606 ), .CO(\mult_x_1/n607 ) );
  CMPR42X1TS \mult_x_1/U412  ( .A(\mult_x_1/n605 ), .B(\mult_x_1/n1006 ), .C(
        \mult_x_1/n615 ), .D(\mult_x_1/n1038 ), .ICI(\mult_x_1/n616 ), .S(
        \mult_x_1/n603 ), .ICO(\mult_x_1/n601 ), .CO(\mult_x_1/n602 ) );
  CMPR42X1TS \mult_x_1/U411  ( .A(\mult_x_1/n603 ), .B(\mult_x_1/n612 ), .C(
        \mult_x_1/n1070 ), .D(\mult_x_1/n1102 ), .ICI(\mult_x_1/n613 ), .S(
        \mult_x_1/n600 ), .ICO(\mult_x_1/n598 ), .CO(\mult_x_1/n599 ) );
  CMPR42X1TS \mult_x_1/U410  ( .A(\mult_x_1/n600 ), .B(\mult_x_1/n609 ), .C(
        \mult_x_1/n1134 ), .D(\mult_x_1/n1166 ), .ICI(\mult_x_1/n610 ), .S(
        \mult_x_1/n597 ), .ICO(\mult_x_1/n595 ), .CO(\mult_x_1/n596 ) );
  CMPR42X1TS \mult_x_1/U409  ( .A(\mult_x_1/n597 ), .B(\mult_x_1/n606 ), .C(
        \mult_x_1/n1198 ), .D(\mult_x_1/n1230 ), .ICI(\mult_x_1/n607 ), .S(
        \mult_x_1/n594 ), .ICO(\mult_x_1/n592 ), .CO(\mult_x_1/n593 ) );
  CMPR42X1TS \mult_x_1/U407  ( .A(\mult_x_1/n591 ), .B(\mult_x_1/n601 ), .C(
        \mult_x_1/n1005 ), .D(\mult_x_1/n1037 ), .ICI(\mult_x_1/n602 ), .S(
        \mult_x_1/n589 ), .ICO(\mult_x_1/n587 ), .CO(\mult_x_1/n588 ) );
  CMPR42X1TS \mult_x_1/U406  ( .A(\mult_x_1/n589 ), .B(\mult_x_1/n598 ), .C(
        \mult_x_1/n1069 ), .D(\mult_x_1/n1101 ), .ICI(\mult_x_1/n599 ), .S(
        \mult_x_1/n586 ), .ICO(\mult_x_1/n584 ), .CO(\mult_x_1/n585 ) );
  CMPR42X1TS \mult_x_1/U405  ( .A(\mult_x_1/n586 ), .B(\mult_x_1/n595 ), .C(
        \mult_x_1/n1133 ), .D(\mult_x_1/n1165 ), .ICI(\mult_x_1/n596 ), .S(
        \mult_x_1/n583 ), .ICO(\mult_x_1/n581 ), .CO(\mult_x_1/n582 ) );
  CMPR42X1TS \mult_x_1/U404  ( .A(\mult_x_1/n583 ), .B(\mult_x_1/n592 ), .C(
        \mult_x_1/n1197 ), .D(\mult_x_1/n1229 ), .ICI(\mult_x_1/n593 ), .S(
        \mult_x_1/n580 ), .ICO(\mult_x_1/n578 ), .CO(\mult_x_1/n579 ) );
  CMPR42X1TS \mult_x_1/U402  ( .A(\mult_x_1/n577 ), .B(\mult_x_1/n587 ), .C(
        \mult_x_1/n1004 ), .D(\mult_x_1/n1036 ), .ICI(\mult_x_1/n588 ), .S(
        \mult_x_1/n575 ), .ICO(\mult_x_1/n573 ), .CO(\mult_x_1/n574 ) );
  CMPR42X1TS \mult_x_1/U401  ( .A(\mult_x_1/n575 ), .B(\mult_x_1/n584 ), .C(
        \mult_x_1/n1068 ), .D(\mult_x_1/n1100 ), .ICI(\mult_x_1/n585 ), .S(
        \mult_x_1/n572 ), .ICO(\mult_x_1/n570 ), .CO(\mult_x_1/n571 ) );
  CMPR42X1TS \mult_x_1/U400  ( .A(\mult_x_1/n572 ), .B(\mult_x_1/n581 ), .C(
        \mult_x_1/n1132 ), .D(\mult_x_1/n1164 ), .ICI(\mult_x_1/n582 ), .S(
        \mult_x_1/n569 ), .ICO(\mult_x_1/n567 ), .CO(\mult_x_1/n568 ) );
  CMPR42X1TS \mult_x_1/U399  ( .A(\mult_x_1/n569 ), .B(\mult_x_1/n578 ), .C(
        \mult_x_1/n1196 ), .D(\mult_x_1/n1228 ), .ICI(\mult_x_1/n579 ), .S(
        \mult_x_1/n566 ), .ICO(\mult_x_1/n564 ), .CO(\mult_x_1/n565 ) );
  CMPR42X1TS \mult_x_1/U397  ( .A(\mult_x_1/n563 ), .B(\mult_x_1/n573 ), .C(
        \mult_x_1/n1003 ), .D(\mult_x_1/n1035 ), .ICI(\mult_x_1/n574 ), .S(
        \mult_x_1/n561 ), .ICO(\mult_x_1/n559 ), .CO(\mult_x_1/n560 ) );
  CMPR42X1TS \mult_x_1/U396  ( .A(\mult_x_1/n561 ), .B(\mult_x_1/n570 ), .C(
        \mult_x_1/n1067 ), .D(\mult_x_1/n1099 ), .ICI(\mult_x_1/n571 ), .S(
        \mult_x_1/n558 ), .ICO(\mult_x_1/n556 ), .CO(\mult_x_1/n557 ) );
  CMPR42X1TS \mult_x_1/U395  ( .A(\mult_x_1/n558 ), .B(\mult_x_1/n567 ), .C(
        \mult_x_1/n1131 ), .D(\mult_x_1/n1163 ), .ICI(\mult_x_1/n568 ), .S(
        \mult_x_1/n555 ), .ICO(\mult_x_1/n553 ), .CO(\mult_x_1/n554 ) );
  CMPR42X1TS \mult_x_1/U394  ( .A(\mult_x_1/n555 ), .B(\mult_x_1/n564 ), .C(
        \mult_x_1/n1195 ), .D(\mult_x_1/n1227 ), .ICI(\mult_x_1/n565 ), .S(
        \mult_x_1/n552 ), .ICO(\mult_x_1/n550 ), .CO(\mult_x_1/n551 ) );
  CMPR42X1TS \mult_x_1/U392  ( .A(\mult_x_1/n549 ), .B(\mult_x_1/n559 ), .C(
        \mult_x_1/n1002 ), .D(\mult_x_1/n1034 ), .ICI(\mult_x_1/n560 ), .S(
        \mult_x_1/n547 ), .ICO(\mult_x_1/n545 ), .CO(\mult_x_1/n546 ) );
  CMPR42X1TS \mult_x_1/U391  ( .A(\mult_x_1/n547 ), .B(\mult_x_1/n556 ), .C(
        \mult_x_1/n1066 ), .D(\mult_x_1/n1098 ), .ICI(\mult_x_1/n557 ), .S(
        \mult_x_1/n544 ), .ICO(\mult_x_1/n542 ), .CO(\mult_x_1/n543 ) );
  CMPR42X1TS \mult_x_1/U390  ( .A(\mult_x_1/n544 ), .B(\mult_x_1/n553 ), .C(
        \mult_x_1/n1130 ), .D(\mult_x_1/n1162 ), .ICI(\mult_x_1/n554 ), .S(
        \mult_x_1/n541 ), .ICO(\mult_x_1/n539 ), .CO(\mult_x_1/n540 ) );
  CMPR42X1TS \mult_x_1/U389  ( .A(\mult_x_1/n541 ), .B(\mult_x_1/n550 ), .C(
        \mult_x_1/n1194 ), .D(\mult_x_1/n1226 ), .ICI(\mult_x_1/n551 ), .S(
        \mult_x_1/n538 ), .ICO(\mult_x_1/n536 ), .CO(\mult_x_1/n537 ) );
  CMPR42X1TS \mult_x_1/U387  ( .A(\mult_x_1/n548 ), .B(\mult_x_1/n535 ), .C(
        \mult_x_1/n545 ), .D(\mult_x_1/n1001 ), .ICI(\mult_x_1/n1033 ), .S(
        \mult_x_1/n533 ), .ICO(\mult_x_1/n531 ), .CO(\mult_x_1/n532 ) );
  CMPR42X1TS \mult_x_1/U386  ( .A(\mult_x_1/n546 ), .B(\mult_x_1/n533 ), .C(
        \mult_x_1/n542 ), .D(\mult_x_1/n1065 ), .ICI(\mult_x_1/n1097 ), .S(
        \mult_x_1/n530 ), .ICO(\mult_x_1/n528 ), .CO(\mult_x_1/n529 ) );
  CMPR42X1TS \mult_x_1/U385  ( .A(\mult_x_1/n543 ), .B(\mult_x_1/n530 ), .C(
        \mult_x_1/n539 ), .D(\mult_x_1/n1129 ), .ICI(\mult_x_1/n1161 ), .S(
        \mult_x_1/n527 ), .ICO(\mult_x_1/n525 ), .CO(\mult_x_1/n526 ) );
  CMPR42X1TS \mult_x_1/U384  ( .A(\mult_x_1/n540 ), .B(\mult_x_1/n527 ), .C(
        \mult_x_1/n536 ), .D(\mult_x_1/n1193 ), .ICI(\mult_x_1/n1225 ), .S(
        \mult_x_1/n524 ), .ICO(\mult_x_1/n522 ), .CO(\mult_x_1/n523 ) );
  CMPR42X1TS \mult_x_1/U382  ( .A(\mult_x_1/n534 ), .B(\mult_x_1/n521 ), .C(
        \mult_x_1/n531 ), .D(\mult_x_1/n1000 ), .ICI(\mult_x_1/n532 ), .S(
        \mult_x_1/n519 ), .ICO(\mult_x_1/n517 ), .CO(\mult_x_1/n518 ) );
  CMPR42X1TS \mult_x_1/U381  ( .A(\mult_x_1/n1032 ), .B(\mult_x_1/n519 ), .C(
        \mult_x_1/n528 ), .D(\mult_x_1/n1064 ), .ICI(\mult_x_1/n529 ), .S(
        \mult_x_1/n516 ), .ICO(\mult_x_1/n514 ), .CO(\mult_x_1/n515 ) );
  CMPR42X1TS \mult_x_1/U380  ( .A(\mult_x_1/n1096 ), .B(\mult_x_1/n516 ), .C(
        \mult_x_1/n525 ), .D(\mult_x_1/n1128 ), .ICI(\mult_x_1/n526 ), .S(
        \mult_x_1/n513 ), .ICO(\mult_x_1/n511 ), .CO(\mult_x_1/n512 ) );
  CMPR42X1TS \mult_x_1/U379  ( .A(\mult_x_1/n1160 ), .B(\mult_x_1/n513 ), .C(
        \mult_x_1/n522 ), .D(\mult_x_1/n1192 ), .ICI(\mult_x_1/n1224 ), .S(
        \mult_x_1/n510 ), .ICO(\mult_x_1/n508 ), .CO(\mult_x_1/n509 ) );
  CMPR42X1TS \mult_x_1/U377  ( .A(\mult_x_1/n520 ), .B(\mult_x_1/n507 ), .C(
        \mult_x_1/n517 ), .D(\mult_x_1/n999 ), .ICI(\mult_x_1/n518 ), .S(
        \mult_x_1/n505 ), .ICO(\mult_x_1/n503 ), .CO(\mult_x_1/n504 ) );
  CMPR42X1TS \mult_x_1/U376  ( .A(\mult_x_1/n1031 ), .B(\mult_x_1/n505 ), .C(
        \mult_x_1/n514 ), .D(\mult_x_1/n1063 ), .ICI(\mult_x_1/n515 ), .S(
        \mult_x_1/n502 ), .ICO(\mult_x_1/n500 ), .CO(\mult_x_1/n501 ) );
  CMPR42X1TS \mult_x_1/U375  ( .A(\mult_x_1/n1095 ), .B(\mult_x_1/n502 ), .C(
        \mult_x_1/n511 ), .D(\mult_x_1/n1127 ), .ICI(\mult_x_1/n512 ), .S(
        \mult_x_1/n499 ), .ICO(\mult_x_1/n497 ), .CO(\mult_x_1/n498 ) );
  CMPR42X1TS \mult_x_1/U374  ( .A(\mult_x_1/n1159 ), .B(\mult_x_1/n499 ), .C(
        \mult_x_1/n508 ), .D(\mult_x_1/n1191 ), .ICI(\mult_x_1/n1223 ), .S(
        \mult_x_1/n496 ), .ICO(\mult_x_1/n494 ), .CO(\mult_x_1/n495 ) );
  CMPR42X1TS \mult_x_1/U372  ( .A(\mult_x_1/n493 ), .B(\mult_x_1/n506 ), .C(
        \mult_x_1/n966 ), .D(\mult_x_1/n503 ), .ICI(\mult_x_1/n998 ), .S(
        \mult_x_1/n491 ), .ICO(\mult_x_1/n489 ), .CO(\mult_x_1/n490 ) );
  CMPR42X1TS \mult_x_1/U371  ( .A(\mult_x_1/n491 ), .B(\mult_x_1/n504 ), .C(
        \mult_x_1/n1030 ), .D(\mult_x_1/n500 ), .ICI(\mult_x_1/n1062 ), .S(
        \mult_x_1/n488 ), .ICO(\mult_x_1/n486 ), .CO(\mult_x_1/n487 ) );
  CMPR42X1TS \mult_x_1/U370  ( .A(\mult_x_1/n488 ), .B(\mult_x_1/n501 ), .C(
        \mult_x_1/n1094 ), .D(\mult_x_1/n497 ), .ICI(\mult_x_1/n1126 ), .S(
        \mult_x_1/n485 ), .ICO(\mult_x_1/n483 ), .CO(\mult_x_1/n484 ) );
  CMPR42X1TS \mult_x_1/U369  ( .A(\mult_x_1/n485 ), .B(\mult_x_1/n498 ), .C(
        \mult_x_1/n1158 ), .D(\mult_x_1/n494 ), .ICI(\mult_x_1/n1190 ), .S(
        \mult_x_1/n482 ), .ICO(\mult_x_1/n480 ), .CO(\mult_x_1/n481 ) );
  CMPR42X1TS \mult_x_1/U367  ( .A(\mult_x_1/n492 ), .B(\mult_x_1/n479 ), .C(
        \mult_x_1/n489 ), .D(\mult_x_1/n965 ), .ICI(\mult_x_1/n490 ), .S(
        \mult_x_1/n478 ), .ICO(\mult_x_1/n476 ), .CO(\mult_x_1/n477 ) );
  CMPR42X1TS \mult_x_1/U366  ( .A(\mult_x_1/n997 ), .B(\mult_x_1/n478 ), .C(
        \mult_x_1/n486 ), .D(\mult_x_1/n1029 ), .ICI(\mult_x_1/n487 ), .S(
        \mult_x_1/n475 ), .ICO(\mult_x_1/n473 ), .CO(\mult_x_1/n474 ) );
  CMPR42X1TS \mult_x_1/U365  ( .A(\mult_x_1/n1061 ), .B(\mult_x_1/n475 ), .C(
        \mult_x_1/n483 ), .D(\mult_x_1/n1093 ), .ICI(\mult_x_1/n484 ), .S(
        \mult_x_1/n472 ), .ICO(\mult_x_1/n470 ), .CO(\mult_x_1/n471 ) );
  CMPR42X1TS \mult_x_1/U364  ( .A(\mult_x_1/n1125 ), .B(\mult_x_1/n472 ), .C(
        \mult_x_1/n480 ), .D(\mult_x_1/n1157 ), .ICI(\mult_x_1/n1189 ), .S(
        \mult_x_1/n469 ), .ICO(\mult_x_1/n467 ), .CO(\mult_x_1/n468 ) );
  CMPR42X1TS \mult_x_1/U362  ( .A(\mult_x_1/n479 ), .B(\mult_x_1/n933 ), .C(
        \mult_x_1/n476 ), .D(\mult_x_1/n964 ), .ICI(\mult_x_1/n477 ), .S(
        \mult_x_1/n464 ), .ICO(\mult_x_1/n462 ), .CO(\mult_x_1/n463 ) );
  CMPR42X1TS \mult_x_1/U361  ( .A(\mult_x_1/n996 ), .B(\mult_x_1/n464 ), .C(
        \mult_x_1/n473 ), .D(\mult_x_1/n1028 ), .ICI(\mult_x_1/n474 ), .S(
        \mult_x_1/n461 ), .ICO(\mult_x_1/n459 ), .CO(\mult_x_1/n460 ) );
  CMPR42X1TS \mult_x_1/U360  ( .A(\mult_x_1/n1060 ), .B(\mult_x_1/n461 ), .C(
        \mult_x_1/n470 ), .D(\mult_x_1/n1092 ), .ICI(\mult_x_1/n471 ), .S(
        \mult_x_1/n458 ), .ICO(\mult_x_1/n456 ), .CO(\mult_x_1/n457 ) );
  CMPR42X1TS \mult_x_1/U359  ( .A(\mult_x_1/n1124 ), .B(\mult_x_1/n458 ), .C(
        \mult_x_1/n467 ), .D(\mult_x_1/n1156 ), .ICI(\mult_x_1/n1188 ), .S(
        \mult_x_1/n455 ), .ICO(\mult_x_1/n453 ), .CO(\mult_x_1/n454 ) );
  CMPR42X1TS \mult_x_1/U358  ( .A(n1674), .B(\mult_x_1/n465 ), .C(
        \mult_x_1/n932 ), .D(\mult_x_1/n462 ), .ICI(\mult_x_1/n963 ), .S(
        \mult_x_1/n452 ), .ICO(\mult_x_1/n428 ), .CO(\mult_x_1/n451 ) );
  CMPR42X1TS \mult_x_1/U357  ( .A(\mult_x_1/n452 ), .B(\mult_x_1/n463 ), .C(
        \mult_x_1/n995 ), .D(\mult_x_1/n459 ), .ICI(\mult_x_1/n1027 ), .S(
        \mult_x_1/n450 ), .ICO(\mult_x_1/n448 ), .CO(\mult_x_1/n449 ) );
  CMPR42X1TS \mult_x_1/U356  ( .A(\mult_x_1/n450 ), .B(\mult_x_1/n460 ), .C(
        \mult_x_1/n1059 ), .D(\mult_x_1/n456 ), .ICI(\mult_x_1/n1091 ), .S(
        \mult_x_1/n447 ), .ICO(\mult_x_1/n445 ), .CO(\mult_x_1/n446 ) );
  CMPR42X1TS \mult_x_1/U355  ( .A(\mult_x_1/n447 ), .B(\mult_x_1/n457 ), .C(
        \mult_x_1/n1123 ), .D(\mult_x_1/n453 ), .ICI(\mult_x_1/n1155 ), .S(
        \mult_x_1/n444 ), .ICO(\mult_x_1/n442 ), .CO(\mult_x_1/n443 ) );
  CMPR42X1TS \mult_x_1/U352  ( .A(\mult_x_1/n451 ), .B(\mult_x_1/n440 ), .C(
        \mult_x_1/n448 ), .D(\mult_x_1/n994 ), .ICI(\mult_x_1/n1026 ), .S(
        \mult_x_1/n438 ), .ICO(\mult_x_1/n436 ), .CO(\mult_x_1/n437 ) );
  CMPR42X1TS \mult_x_1/U351  ( .A(\mult_x_1/n449 ), .B(\mult_x_1/n438 ), .C(
        \mult_x_1/n445 ), .D(\mult_x_1/n1058 ), .ICI(\mult_x_1/n1090 ), .S(
        \mult_x_1/n435 ), .ICO(\mult_x_1/n433 ), .CO(\mult_x_1/n434 ) );
  CMPR42X1TS \mult_x_1/U350  ( .A(\mult_x_1/n446 ), .B(\mult_x_1/n435 ), .C(
        \mult_x_1/n442 ), .D(\mult_x_1/n1122 ), .ICI(\mult_x_1/n1154 ), .S(
        \mult_x_1/n432 ), .ICO(\mult_x_1/n430 ), .CO(\mult_x_1/n431 ) );
  CMPR42X1TS \mult_x_1/U347  ( .A(\mult_x_1/n439 ), .B(\mult_x_1/n427 ), .C(
        \mult_x_1/n436 ), .D(\mult_x_1/n993 ), .ICI(\mult_x_1/n437 ), .S(
        \mult_x_1/n425 ), .ICO(\mult_x_1/n423 ), .CO(\mult_x_1/n424 ) );
  CMPR42X1TS \mult_x_1/U346  ( .A(\mult_x_1/n1025 ), .B(\mult_x_1/n425 ), .C(
        \mult_x_1/n433 ), .D(\mult_x_1/n1057 ), .ICI(\mult_x_1/n434 ), .S(
        \mult_x_1/n422 ), .ICO(\mult_x_1/n420 ), .CO(\mult_x_1/n421 ) );
  CMPR42X1TS \mult_x_1/U345  ( .A(\mult_x_1/n1089 ), .B(\mult_x_1/n422 ), .C(
        \mult_x_1/n430 ), .D(\mult_x_1/n1121 ), .ICI(\mult_x_1/n1153 ), .S(
        \mult_x_1/n419 ), .ICO(\mult_x_1/n417 ), .CO(\mult_x_1/n418 ) );
  CMPR42X1TS \mult_x_1/U343  ( .A(\mult_x_1/n416 ), .B(\mult_x_1/n960 ), .C(
        \mult_x_1/n426 ), .D(\mult_x_1/n423 ), .ICI(\mult_x_1/n992 ), .S(
        \mult_x_1/n414 ), .ICO(\mult_x_1/n412 ), .CO(\mult_x_1/n413 ) );
  CMPR42X1TS \mult_x_1/U342  ( .A(\mult_x_1/n414 ), .B(\mult_x_1/n424 ), .C(
        \mult_x_1/n1024 ), .D(\mult_x_1/n420 ), .ICI(\mult_x_1/n1056 ), .S(
        \mult_x_1/n411 ), .ICO(\mult_x_1/n409 ), .CO(\mult_x_1/n410 ) );
  CMPR42X1TS \mult_x_1/U341  ( .A(\mult_x_1/n411 ), .B(\mult_x_1/n421 ), .C(
        \mult_x_1/n1088 ), .D(\mult_x_1/n417 ), .ICI(\mult_x_1/n1120 ), .S(
        \mult_x_1/n408 ), .ICO(\mult_x_1/n406 ), .CO(\mult_x_1/n407 ) );
  CMPR42X1TS \mult_x_1/U339  ( .A(\mult_x_1/n415 ), .B(\mult_x_1/n405 ), .C(
        \mult_x_1/n412 ), .D(\mult_x_1/n959 ), .ICI(\mult_x_1/n991 ), .S(
        \mult_x_1/n404 ), .ICO(\mult_x_1/n402 ), .CO(\mult_x_1/n403 ) );
  CMPR42X1TS \mult_x_1/U338  ( .A(\mult_x_1/n413 ), .B(\mult_x_1/n404 ), .C(
        \mult_x_1/n409 ), .D(\mult_x_1/n1023 ), .ICI(\mult_x_1/n1055 ), .S(
        \mult_x_1/n401 ), .ICO(\mult_x_1/n399 ), .CO(\mult_x_1/n400 ) );
  CMPR42X1TS \mult_x_1/U337  ( .A(\mult_x_1/n410 ), .B(\mult_x_1/n401 ), .C(
        \mult_x_1/n406 ), .D(\mult_x_1/n1087 ), .ICI(\mult_x_1/n1119 ), .S(
        \mult_x_1/n398 ), .ICO(\mult_x_1/n396 ), .CO(\mult_x_1/n397 ) );
  CMPR42X1TS \mult_x_1/U335  ( .A(\mult_x_1/n405 ), .B(\mult_x_1/n928 ), .C(
        \mult_x_1/n402 ), .D(\mult_x_1/n958 ), .ICI(\mult_x_1/n403 ), .S(
        \mult_x_1/n393 ), .ICO(\mult_x_1/n391 ), .CO(\mult_x_1/n392 ) );
  CMPR42X1TS \mult_x_1/U334  ( .A(\mult_x_1/n990 ), .B(\mult_x_1/n393 ), .C(
        \mult_x_1/n399 ), .D(\mult_x_1/n1022 ), .ICI(\mult_x_1/n400 ), .S(
        \mult_x_1/n390 ), .ICO(\mult_x_1/n388 ), .CO(\mult_x_1/n389 ) );
  CMPR42X1TS \mult_x_1/U333  ( .A(\mult_x_1/n1054 ), .B(\mult_x_1/n390 ), .C(
        \mult_x_1/n396 ), .D(\mult_x_1/n1086 ), .ICI(\mult_x_1/n1118 ), .S(
        \mult_x_1/n387 ), .ICO(\mult_x_1/n385 ), .CO(\mult_x_1/n386 ) );
  CMPR42X1TS \mult_x_1/U332  ( .A(n1673), .B(\mult_x_1/n394 ), .C(
        \mult_x_1/n927 ), .D(\mult_x_1/n391 ), .ICI(\mult_x_1/n957 ), .S(
        \mult_x_1/n384 ), .ICO(\mult_x_1/n366 ), .CO(\mult_x_1/n383 ) );
  CMPR42X1TS \mult_x_1/U331  ( .A(\mult_x_1/n384 ), .B(\mult_x_1/n392 ), .C(
        \mult_x_1/n989 ), .D(\mult_x_1/n388 ), .ICI(\mult_x_1/n1021 ), .S(
        \mult_x_1/n382 ), .ICO(\mult_x_1/n380 ), .CO(\mult_x_1/n381 ) );
  CMPR42X1TS \mult_x_1/U330  ( .A(\mult_x_1/n382 ), .B(\mult_x_1/n389 ), .C(
        \mult_x_1/n1053 ), .D(\mult_x_1/n385 ), .ICI(\mult_x_1/n1085 ), .S(
        \mult_x_1/n379 ), .ICO(\mult_x_1/n377 ), .CO(\mult_x_1/n378 ) );
  CMPR42X1TS \mult_x_1/U327  ( .A(\mult_x_1/n383 ), .B(\mult_x_1/n375 ), .C(
        \mult_x_1/n380 ), .D(\mult_x_1/n988 ), .ICI(\mult_x_1/n1020 ), .S(
        \mult_x_1/n373 ), .ICO(\mult_x_1/n371 ), .CO(\mult_x_1/n372 ) );
  CMPR42X1TS \mult_x_1/U326  ( .A(\mult_x_1/n381 ), .B(\mult_x_1/n373 ), .C(
        \mult_x_1/n377 ), .D(\mult_x_1/n1052 ), .ICI(\mult_x_1/n1084 ), .S(
        \mult_x_1/n370 ), .ICO(\mult_x_1/n368 ), .CO(\mult_x_1/n369 ) );
  CMPR42X1TS \mult_x_1/U323  ( .A(\mult_x_1/n374 ), .B(\mult_x_1/n365 ), .C(
        \mult_x_1/n371 ), .D(\mult_x_1/n987 ), .ICI(\mult_x_1/n372 ), .S(
        \mult_x_1/n363 ), .ICO(\mult_x_1/n361 ), .CO(\mult_x_1/n362 ) );
  CMPR42X1TS \mult_x_1/U322  ( .A(\mult_x_1/n1019 ), .B(\mult_x_1/n363 ), .C(
        \mult_x_1/n368 ), .D(\mult_x_1/n1051 ), .ICI(\mult_x_1/n1083 ), .S(
        \mult_x_1/n360 ), .ICO(\mult_x_1/n358 ), .CO(\mult_x_1/n359 ) );
  CMPR42X1TS \mult_x_1/U320  ( .A(\mult_x_1/n357 ), .B(\mult_x_1/n364 ), .C(
        \mult_x_1/n954 ), .D(\mult_x_1/n361 ), .ICI(\mult_x_1/n986 ), .S(
        \mult_x_1/n355 ), .ICO(\mult_x_1/n353 ), .CO(\mult_x_1/n354 ) );
  CMPR42X1TS \mult_x_1/U319  ( .A(\mult_x_1/n355 ), .B(\mult_x_1/n362 ), .C(
        \mult_x_1/n1018 ), .D(\mult_x_1/n358 ), .ICI(\mult_x_1/n1050 ), .S(
        \mult_x_1/n352 ), .ICO(\mult_x_1/n350 ), .CO(\mult_x_1/n351 ) );
  CMPR42X1TS \mult_x_1/U317  ( .A(\mult_x_1/n356 ), .B(\mult_x_1/n349 ), .C(
        \mult_x_1/n353 ), .D(\mult_x_1/n953 ), .ICI(\mult_x_1/n985 ), .S(
        \mult_x_1/n348 ), .ICO(\mult_x_1/n346 ), .CO(\mult_x_1/n347 ) );
  CMPR42X1TS \mult_x_1/U316  ( .A(\mult_x_1/n354 ), .B(\mult_x_1/n348 ), .C(
        \mult_x_1/n350 ), .D(\mult_x_1/n1017 ), .ICI(\mult_x_1/n1049 ), .S(
        \mult_x_1/n345 ), .ICO(\mult_x_1/n343 ), .CO(\mult_x_1/n344 ) );
  CMPR42X1TS \mult_x_1/U314  ( .A(\mult_x_1/n349 ), .B(\mult_x_1/n923 ), .C(
        \mult_x_1/n346 ), .D(\mult_x_1/n952 ), .ICI(\mult_x_1/n347 ), .S(
        \mult_x_1/n340 ), .ICO(\mult_x_1/n338 ), .CO(\mult_x_1/n339 ) );
  CMPR42X1TS \mult_x_1/U313  ( .A(\mult_x_1/n984 ), .B(\mult_x_1/n340 ), .C(
        \mult_x_1/n343 ), .D(\mult_x_1/n1016 ), .ICI(\mult_x_1/n1048 ), .S(
        \mult_x_1/n337 ), .ICO(\mult_x_1/n335 ), .CO(\mult_x_1/n336 ) );
  CMPR42X1TS \mult_x_1/U312  ( .A(n1672), .B(\mult_x_1/n341 ), .C(
        \mult_x_1/n922 ), .D(\mult_x_1/n338 ), .ICI(\mult_x_1/n951 ), .S(
        \mult_x_1/n334 ), .ICO(\mult_x_1/n322 ), .CO(\mult_x_1/n333 ) );
  CMPR42X1TS \mult_x_1/U311  ( .A(\mult_x_1/n334 ), .B(\mult_x_1/n339 ), .C(
        \mult_x_1/n983 ), .D(\mult_x_1/n335 ), .ICI(\mult_x_1/n1015 ), .S(
        \mult_x_1/n332 ), .ICO(\mult_x_1/n330 ), .CO(\mult_x_1/n331 ) );
  CMPR42X1TS \mult_x_1/U308  ( .A(\mult_x_1/n333 ), .B(\mult_x_1/n328 ), .C(
        \mult_x_1/n330 ), .D(\mult_x_1/n982 ), .ICI(\mult_x_1/n1014 ), .S(
        \mult_x_1/n326 ), .ICO(\mult_x_1/n324 ), .CO(\mult_x_1/n325 ) );
  CMPR42X1TS \mult_x_1/U305  ( .A(\mult_x_1/n949 ), .B(\mult_x_1/n321 ), .C(
        \mult_x_1/n324 ), .D(\mult_x_1/n981 ), .ICI(\mult_x_1/n1013 ), .S(
        \mult_x_1/n319 ), .ICO(\mult_x_1/n317 ), .CO(\mult_x_1/n318 ) );
  CMPR42X1TS \mult_x_1/U303  ( .A(\mult_x_1/n316 ), .B(\mult_x_1/n320 ), .C(
        \mult_x_1/n948 ), .D(\mult_x_1/n317 ), .ICI(\mult_x_1/n980 ), .S(
        \mult_x_1/n315 ), .ICO(\mult_x_1/n313 ), .CO(\mult_x_1/n314 ) );
  CMPR42X1TS \mult_x_1/U301  ( .A(\mult_x_1/n918 ), .B(\mult_x_1/n312 ), .C(
        \mult_x_1/n313 ), .D(\mult_x_1/n947 ), .ICI(\mult_x_1/n979 ), .S(
        \mult_x_1/n311 ), .ICO(\mult_x_1/n309 ), .CO(\mult_x_1/n310 ) );
  CMPR42X1TS \mult_x_1/U299  ( .A(\mult_x_1/n312 ), .B(\mult_x_1/n917 ), .C(
        \mult_x_1/n309 ), .D(\mult_x_1/n946 ), .ICI(\mult_x_1/n978 ), .S(
        \mult_x_1/n306 ), .ICO(\mult_x_1/n304 ), .CO(\mult_x_1/n305 ) );
  CMPR42X1TS \mult_x_1/U298  ( .A(n1671), .B(\mult_x_1/n307 ), .C(
        \mult_x_1/n916 ), .D(\mult_x_1/n304 ), .ICI(\mult_x_1/n945 ), .S(
        \mult_x_1/n303 ), .ICO(\mult_x_1/n297 ), .CO(\mult_x_1/n302 ) );
  CMPR32X2TS U1 ( .A(n1375), .B(n1374), .C(n1373), .CO(n1389), .S(n1345) );
  CMPR32X2TS U2 ( .A(B[13]), .B(B[14]), .C(n166), .CO(n175), .S(n158) );
  CMPR32X2TS U3 ( .A(n1551), .B(n1550), .C(n1549), .CO(n1574), .S(n1544) );
  CLKAND2X2TS U4 ( .A(n985), .B(n543), .Y(n540) );
  NAND2BX2TS U5 ( .AN(n499), .B(n1012), .Y(n1643) );
  NAND2BX2TS U6 ( .AN(n998), .B(n1515), .Y(n1652) );
  CLKAND2X2TS U7 ( .A(A[0]), .B(n5), .Y(n2) );
  NAND2BX2TS U8 ( .AN(n999), .B(n997), .Y(n1518) );
  CLKAND2X2TS U9 ( .A(n18), .B(n19), .Y(n15) );
  NAND2X2TS U10 ( .A(n94), .B(n95), .Y(n1279) );
  NAND2X2TS U11 ( .A(n719), .B(n718), .Y(n1264) );
  NAND2X2TS U12 ( .A(n500), .B(n498), .Y(n723) );
  NAND2X2TS U13 ( .A(n321), .B(n320), .Y(n322) );
  NAND2BX2TS U14 ( .AN(n500), .B(n498), .Y(n727) );
  CLKAND2X2TS U15 ( .A(A[1]), .B(n8), .Y(n4) );
  NAND3X2TS U16 ( .A(A[29]), .B(A[30]), .C(A[31]), .Y(n1559) );
  INVX3TS U17 ( .A(A[20]), .Y(n1672) );
  CLKINVX3TS U18 ( .A(A[17]), .Y(n539) );
  INVX3TS U19 ( .A(A[14]), .Y(n1673) );
  CLKINVX3TS U20 ( .A(A[11]), .Y(n1638) );
  CLKINVX3TS U21 ( .A(A[8]), .Y(n1674) );
  CLKINVX3TS U22 ( .A(A[23]), .Y(n1621) );
  INVX3TS U23 ( .A(A[26]), .Y(n1671) );
  CLKINVX3TS U24 ( .A(A[5]), .Y(n14) );
  ADDFX1TS U25 ( .A(n1033), .B(n1032), .CI(n1031), .CO(n1085), .S(n1022) );
  ADDFX1TS U26 ( .A(n843), .B(n842), .CI(n841), .CO(n845), .S(n844) );
  ADDFX1TS U27 ( .A(n847), .B(n846), .CI(n845), .CO(n834), .S(n848) );
  ADDFX1TS U28 ( .A(n836), .B(n835), .CI(n834), .CO(n800), .S(n837) );
  ADDFX1TS U29 ( .A(n693), .B(n692), .CI(n691), .CO(n662), .S(n694) );
  ADDFX1TS U30 ( .A(n693), .B(n689), .CI(n688), .CO(n648), .S(n690) );
  ADDFX1TS U31 ( .A(n693), .B(n686), .CI(n685), .CO(n668), .S(n687) );
  ADDFX1TS U32 ( .A(A[5]), .B(A[2]), .CI(n571), .CO(n514), .S(n572) );
  ADDFX1TS U33 ( .A(n1086), .B(n1085), .CI(n1084), .CO(n1037), .S(n1087) );
  ADDFX1TS U34 ( .A(\mult_x_1/n428 ), .B(n586), .CI(n585), .CO(n563), .S(n587)
         );
  ADDFX1TS U35 ( .A(\mult_x_1/n428 ), .B(n589), .CI(n588), .CO(n554), .S(n590)
         );
  ADDFX1TS U36 ( .A(A[11]), .B(n471), .CI(n470), .CO(n417), .S(n472) );
  ADDFX1TS U37 ( .A(B[24]), .B(B[25]), .CI(n263), .CO(n258), .S(n264) );
  ADDFX1TS U38 ( .A(B[3]), .B(B[4]), .CI(n46), .CO(n58), .S(n31) );
  ADDFX1TS U39 ( .A(B[4]), .B(B[5]), .CI(n58), .CO(n79), .S(n47) );
  ADDFX1TS U40 ( .A(B[5]), .B(B[6]), .CI(n79), .CO(n88), .S(n59) );
  ADDFX1TS U41 ( .A(B[6]), .B(B[7]), .CI(n88), .CO(n111), .S(n80) );
  ADDFX1TS U42 ( .A(B[7]), .B(B[8]), .CI(n111), .CO(n117), .S(n89) );
  ADDFX1TS U43 ( .A(B[9]), .B(B[10]), .CI(n130), .CO(n139), .S(n112) );
  ADDFX1TS U44 ( .A(B[10]), .B(B[11]), .CI(n139), .CO(n148), .S(n131) );
  ADDFX1TS U45 ( .A(B[12]), .B(B[13]), .CI(n157), .CO(n166), .S(n149) );
  ADDFX1TS U46 ( .A(B[11]), .B(B[12]), .CI(n148), .CO(n157), .S(n140) );
  ADDFX1TS U47 ( .A(B[15]), .B(B[16]), .CI(n184), .CO(n193), .S(n176) );
  ADDFX1TS U48 ( .A(B[14]), .B(B[15]), .CI(n175), .CO(n184), .S(n167) );
  ADDFX1TS U49 ( .A(B[16]), .B(B[17]), .CI(n193), .CO(n202), .S(n185) );
  ADDFX1TS U50 ( .A(n1360), .B(n1359), .CI(n1358), .CO(n1367), .S(n1353) );
  ADDFX1TS U51 ( .A(B[18]), .B(B[19]), .CI(n211), .CO(n220), .S(n203) );
  ADDFX1TS U52 ( .A(B[17]), .B(B[18]), .CI(n202), .CO(n211), .S(n194) );
  ADDFX1TS U53 ( .A(n1368), .B(n1367), .CI(n1366), .CO(n1365), .S(n1369) );
  ADDFX1TS U54 ( .A(B[19]), .B(B[20]), .CI(n220), .CO(n229), .S(n212) );
  ADDFX1TS U55 ( .A(B[20]), .B(B[21]), .CI(n229), .CO(n278), .S(n221) );
  ADDFX1TS U56 ( .A(B[21]), .B(B[22]), .CI(n278), .CO(n273), .S(n279) );
  ADDFX1TS U57 ( .A(B[22]), .B(B[23]), .CI(n273), .CO(n268), .S(n274) );
  ADDFX1TS U58 ( .A(B[23]), .B(B[24]), .CI(n268), .CO(n263), .S(n269) );
  ADDFX1TS U59 ( .A(B[25]), .B(B[26]), .CI(n258), .CO(n253), .S(n259) );
  ADDFX1TS U60 ( .A(B[26]), .B(B[27]), .CI(n253), .CO(n248), .S(n254) );
  ADDFX1TS U61 ( .A(B[27]), .B(B[28]), .CI(n248), .CO(n243), .S(n249) );
  ADDFX1TS U62 ( .A(B[28]), .B(B[29]), .CI(n243), .CO(n238), .S(n244) );
  ADDFX1TS U63 ( .A(\mult_x_1/n366 ), .B(n487), .CI(n486), .CO(n465), .S(n488)
         );
  ADDFX1TS U64 ( .A(\mult_x_1/n366 ), .B(n490), .CI(n489), .CO(n455), .S(n491)
         );
  ADDFX1TS U65 ( .A(A[17]), .B(n372), .CI(n371), .CO(n346), .S(n373) );
  ADDFX1TS U66 ( .A(B[8]), .B(B[9]), .CI(n117), .CO(n130), .S(n118) );
  ADDFX1TS U67 ( .A(B[2]), .B(B[3]), .CI(n30), .CO(n46), .S(n22) );
  ADDFX1TS U68 ( .A(n1575), .B(n1574), .CI(n1573), .CO(n1558), .S(n1576) );
  ADDFX1TS U69 ( .A(B[29]), .B(B[30]), .CI(n238), .CO(n233), .S(n239) );
  ADDFX1TS U70 ( .A(\mult_x_1/n322 ), .B(n399), .CI(n398), .CO(n419), .S(n400)
         );
  ADDFX1TS U71 ( .A(\mult_x_1/n322 ), .B(n419), .CI(n418), .CO(n381), .S(n420)
         );
  ADDFX1TS U72 ( .A(n1621), .B(\mult_x_1/n322 ), .CI(n1620), .CO(
        \mult_x_1/n307 ), .S(\mult_x_1/n316 ) );
  ADDFX1TS U73 ( .A(n103), .B(n102), .CI(n101), .CO(n1598), .S(n109) );
  ADDFX1TS U74 ( .A(n1599), .B(n1598), .CI(n1597), .CO(n1600), .S(n123) );
  ADDFX1TS U75 ( .A(n365), .B(n364), .CI(n363), .CO(n350), .S(n366) );
  ADDFX1TS U76 ( .A(B[30]), .B(B[31]), .CI(n233), .CO(n230), .S(n234) );
  ADDFX1TS U77 ( .A(\mult_x_1/n297 ), .B(n1568), .CI(n1567), .CO(n1586), .S(
        n1570) );
  ADDFX1TS U78 ( .A(\mult_x_1/n297 ), .B(n1578), .CI(n1577), .CO(n1595), .S(
        n1587) );
  ADDFX1TS U79 ( .A(A[29]), .B(n1590), .CI(n1589), .CO(n1666), .S(n1594) );
  ADDFX1TS U80 ( .A(n52), .B(n1613), .CI(n51), .CO(n63), .S(n35) );
  ADDFX1TS U81 ( .A(n65), .B(n64), .CI(n63), .CO(n84), .S(n53) );
  ADDFX1TS U82 ( .A(n86), .B(n85), .CI(n84), .CO(n107), .S(n66) );
  ADDFX1TS U83 ( .A(n109), .B(n108), .CI(n107), .CO(n122), .S(n87) );
  ADDFX1TS U84 ( .A(n124), .B(n123), .CI(n122), .CO(n126), .S(n110) );
  ADDFX1TS U85 ( .A(n137), .B(n136), .CI(n135), .CO(n144), .S(n125) );
  ADDFX1TS U86 ( .A(n146), .B(n145), .CI(n144), .CO(n153), .S(n138) );
  ADDFX1TS U87 ( .A(n164), .B(n163), .CI(n162), .CO(n171), .S(n156) );
  ADDFX1TS U88 ( .A(n155), .B(n154), .CI(n153), .CO(n162), .S(n147) );
  ADDFX1TS U89 ( .A(n191), .B(n190), .CI(n189), .CO(n198), .S(n183) );
  ADDFX1TS U90 ( .A(n173), .B(n172), .CI(n171), .CO(n180), .S(n165) );
  ADDFX1TS U91 ( .A(n182), .B(n181), .CI(n180), .CO(n189), .S(n174) );
  ADDFX1TS U92 ( .A(n200), .B(n199), .CI(n198), .CO(n207), .S(n192) );
  ADDFX1TS U93 ( .A(n218), .B(n217), .CI(n216), .CO(n225), .S(n210) );
  ADDFX1TS U94 ( .A(n209), .B(n208), .CI(n207), .CO(n216), .S(n201) );
  ADDFX1TS U95 ( .A(n227), .B(n226), .CI(n225), .CO(n285), .S(n219) );
  ADDFX1TS U96 ( .A(n287), .B(n286), .CI(n285), .CO(n306), .S(n228) );
  ADDFX1TS U97 ( .A(n308), .B(n307), .CI(n306), .CO(n314), .S(n309) );
  ADDFX1TS U98 ( .A(n316), .B(n315), .CI(n314), .CO(n334), .S(n317) );
  ADDFX1TS U99 ( .A(n336), .B(n335), .CI(n334), .CO(n363), .S(n337) );
  ADDFX1TS U100 ( .A(n352), .B(n351), .CI(n350), .CO(n367), .S(n353) );
  ADDFX1TS U101 ( .A(n369), .B(n368), .CI(n367), .CO(n439), .S(n370) );
  ADDFX1TS U102 ( .A(n441), .B(n440), .CI(n439), .CO(n446), .S(n442) );
  ADDFX1TS U103 ( .A(n448), .B(n447), .CI(n446), .CO(n456), .S(n449) );
  ADDFX1TS U104 ( .A(n458), .B(n457), .CI(n456), .CO(n494), .S(n459) );
  ADDFX1TS U105 ( .A(n496), .B(n495), .CI(n494), .CO(n302), .S(n497) );
  ADDFX1TS U106 ( .A(n1070), .B(n1069), .CI(n1068), .CO(n1157), .S(n996) );
  ADDFX1TS U107 ( .A(n1344), .B(n1343), .CI(n1342), .CO(n1373), .S(n1259) );
  ADDFX1TS U108 ( .A(n677), .B(n676), .CI(n675), .CO(n713), .S(n652) );
  ADDFX1TS U109 ( .A(n974), .B(n973), .CI(n972), .CO(n993), .S(n952) );
  ADDFX1TS U110 ( .A(n832), .B(n831), .CI(n830), .CO(n949), .S(n820) );
  ADDFX1TS U111 ( .A(n1587), .B(n1586), .CI(n1585), .CO(n1593), .S(n1572) );
  ADDFX1TS U112 ( .A(n739), .B(n738), .CI(n737), .CO(n817), .S(n716) );
  ADDFX1TS U113 ( .A(n1170), .B(n1169), .CI(n1168), .CO(n1256), .S(n1160) );
  ADDFX1TS U114 ( .A(n1391), .B(n1390), .CI(n1389), .CO(n1569), .S(n1376) );
  ADDFX1TS U115 ( .A(n1666), .B(n1667), .CI(n1665), .CO(n1668), .S(n1596) );
  ADDFX1TS U116 ( .A(n304), .B(n303), .CI(n302), .CO(n310), .S(n288) );
  ADDFX1TS U117 ( .A(n569), .B(n568), .CI(n567), .CO(n594), .S(n518) );
  ADDFX1TS U118 ( .A(n484), .B(n483), .CI(n482), .CO(n515), .S(n469) );
  ADDFX1TS U119 ( .A(n312), .B(n311), .CI(n310), .CO(n330), .S(n305) );
  ADDFX1TS U120 ( .A(n596), .B(n595), .CI(n594), .CO(n649), .S(n570) );
  ADDFX1TS U121 ( .A(n407), .B(n406), .CI(n405), .CO(n466), .S(n388) );
  ADDFX1TS U122 ( .A(n361), .B(n360), .CI(n359), .CO(n385), .S(n333) );
  ADDFX1TS U123 ( .A(n332), .B(n331), .CI(n330), .CO(n359), .S(n313) );
  ADDFX1TS U124 ( .A(n387), .B(n386), .CI(n385), .CO(n405), .S(n362) );
  ADDFX1TS U125 ( .A(n468), .B(n467), .CI(n466), .CO(n482), .S(n408) );
  ADDFX1TS U126 ( .A(n651), .B(n650), .CI(n649), .CO(n675), .S(n597) );
  ADDFX1TS U127 ( .A(n715), .B(n714), .CI(n713), .CO(n737), .S(n678) );
  ADDFX1TS U128 ( .A(n819), .B(n818), .CI(n817), .CO(n830), .S(n740) );
  ADDFX1TS U129 ( .A(n951), .B(n950), .CI(n949), .CO(n972), .S(n833) );
  ADDFX1TS U130 ( .A(n995), .B(n994), .CI(n993), .CO(n1068), .S(n975) );
  ADDFX1TS U131 ( .A(n1159), .B(n1158), .CI(n1157), .CO(n1168), .S(n1071) );
  ADDFX1TS U132 ( .A(n1258), .B(n1257), .CI(n1256), .CO(n1342), .S(n1171) );
  ADDFX1TS U133 ( .A(n1571), .B(n1570), .CI(n1569), .CO(n1585), .S(n1392) );
  ADDFX1TS U134 ( .A(n1595), .B(n1594), .CI(n1593), .CO(n1665), .S(n1588) );
  ADDFX1TS U135 ( .A(n517), .B(n516), .CI(n515), .CO(n567), .S(n485) );
  ADDFX1TS U136 ( .A(n128), .B(n127), .CI(n126), .CO(n135), .S(n129) );
  AND3X1TS U137 ( .A(n857), .B(n771), .C(n770), .Y(n1) );
  INVX2TS U138 ( .A(A[2]), .Y(n693) );
  INVX2TS U139 ( .A(n693), .Y(n1616) );
  AOI2BB2XLTS U140 ( .B0(n1616), .B1(A[1]), .A0N(A[1]), .A1N(n1616), .Y(n5) );
  INVX2TS U141 ( .A(n2), .Y(n300) );
  INVX2TS U142 ( .A(B[2]), .Y(n29) );
  INVX2TS U143 ( .A(B[1]), .Y(n23) );
  OAI21XLTS U144 ( .A0(B[0]), .A1(n23), .B0(n29), .Y(n3) );
  OAI31X2TS U145 ( .A0(B[0]), .A1(n29), .A2(n23), .B0(n3), .Y(n1517) );
  INVX2TS U146 ( .A(A[0]), .Y(n8) );
  NOR3XLTS U147 ( .A(A[0]), .B(A[1]), .C(n693), .Y(n231) );
  AOI22X1TS U148 ( .A0(n4), .A1(B[1]), .B0(n231), .B1(B[0]), .Y(n7) );
  NOR2XLTS U149 ( .A(n8), .B(n5), .Y(n24) );
  NAND2X1TS U150 ( .A(n24), .B(B[2]), .Y(n6) );
  OAI211XLTS U151 ( .A0(n300), .A1(n1517), .B0(n7), .C0(n6), .Y(n13) );
  INVX2TS U152 ( .A(B[0]), .Y(n9) );
  NOR2XLTS U153 ( .A(n8), .B(n9), .Y(Product[0]) );
  OAI22X1TS U154 ( .A0(n23), .A1(n9), .B0(B[0]), .B1(B[1]), .Y(n1516) );
  INVX2TS U155 ( .A(n1516), .Y(n1183) );
  AOI222XLTS U156 ( .A0(n24), .A1(B[1]), .B0(n4), .B1(B[0]), .C0(n2), .C1(
        n1183), .Y(n1619) );
  OAI2BB1X1TS U157 ( .A0N(n1616), .A1N(Product[0]), .B0(n1619), .Y(n1617) );
  NOR2XLTS U158 ( .A(n693), .B(n1617), .Y(n11) );
  INVX2TS U159 ( .A(n13), .Y(n10) );
  NAND2X1TS U160 ( .A(n11), .B(n10), .Y(n28) );
  OAI21XLTS U161 ( .A0(n13), .A1(n1616), .B0(n28), .Y(n12) );
  AOI31XLTS U162 ( .A0(n13), .A1(n1616), .A2(n1617), .B0(n12), .Y(Product[2])
         );
  INVX2TS U163 ( .A(A[4]), .Y(n17) );
  OAI22X1TS U164 ( .A0(n14), .A1(n17), .B0(A[4]), .B1(A[5]), .Y(n18) );
  INVX2TS U165 ( .A(A[3]), .Y(n16) );
  OAI22X1TS U166 ( .A0(n693), .A1(A[3]), .B0(n16), .B1(n1616), .Y(n19) );
  AOI22X1TS U167 ( .A0(A[3]), .A1(n17), .B0(A[4]), .B1(n16), .Y(n36) );
  NOR2XLTS U168 ( .A(n19), .B(n36), .Y(n1512) );
  INVX2TS U169 ( .A(n18), .Y(n38) );
  CLKAND2X2TS U170 ( .A(n19), .B(n38), .Y(n1513) );
  AOI222XLTS U171 ( .A0(B[1]), .A1(n15), .B0(B[0]), .B1(n1512), .C0(n1183), 
        .C1(n1513), .Y(n21) );
  NAND3XLTS U172 ( .A(B[0]), .B(n19), .C(A[5]), .Y(n20) );
  INVX2TS U173 ( .A(n19), .Y(n37) );
  OAI31X1TS U174 ( .A0(n9), .A1(n37), .A2(n14), .B0(n21), .Y(n43) );
  OAI21XLTS U175 ( .A0(n21), .A1(n20), .B0(n43), .Y(n52) );
  AOI21X1TS U176 ( .A0(n29), .A1(n9), .B0(n23), .Y(n30) );
  INVX2TS U177 ( .A(n22), .Y(n1527) );
  INVX2TS U178 ( .A(n231), .Y(n113) );
  OAI22X1TS U179 ( .A0(n1527), .A1(n300), .B0(n23), .B1(n113), .Y(n27) );
  INVX2TS U180 ( .A(B[3]), .Y(n1554) );
  INVX2TS U181 ( .A(n24), .Y(n281) );
  INVX2TS U182 ( .A(n4), .Y(n280) );
  OAI22X1TS U183 ( .A0(n1554), .A1(n281), .B0(n29), .B1(n280), .Y(n26) );
  OAI21XLTS U184 ( .A0(n27), .A1(n26), .B0(n693), .Y(n25) );
  OAI31X1TS U185 ( .A0(n27), .A1(n693), .A2(n26), .B0(n25), .Y(n1614) );
  OAI21XLTS U186 ( .A0(n9), .A1(n37), .B0(n28), .Y(n1615) );
  NAND2X1TS U187 ( .A(n1614), .B(n1615), .Y(n1613) );
  INVX2TS U188 ( .A(n31), .Y(n1537) );
  OAI22X1TS U189 ( .A0(n29), .A1(n113), .B0(n300), .B1(n1537), .Y(n34) );
  INVX2TS U190 ( .A(B[4]), .Y(n813) );
  OAI22X1TS U191 ( .A0(n1554), .A1(n280), .B0(n281), .B1(n813), .Y(n33) );
  OAI21XLTS U192 ( .A0(n34), .A1(n33), .B0(n1616), .Y(n32) );
  OAI31X1TS U193 ( .A0(n34), .A1(n1616), .A2(n33), .B0(n32), .Y(n51) );
  INVX2TS U194 ( .A(n35), .Y(Product[4]) );
  INVX2TS U195 ( .A(n1512), .Y(n1496) );
  AND3X1TS U196 ( .A(n38), .B(n37), .C(n36), .Y(n1511) );
  INVX2TS U197 ( .A(n1511), .Y(n1659) );
  INVX2TS U198 ( .A(n1513), .Y(n1660) );
  OAI22X1TS U199 ( .A0(n9), .A1(n1659), .B0(n1517), .B1(n1660), .Y(n39) );
  AOI21X1TS U200 ( .A0(B[2]), .A1(n15), .B0(n39), .Y(n40) );
  OAI21XLTS U201 ( .A0(n23), .A1(n1496), .B0(n40), .Y(n45) );
  NOR2XLTS U202 ( .A(n14), .B(n43), .Y(n42) );
  INVX2TS U203 ( .A(n45), .Y(n41) );
  NAND2X1TS U204 ( .A(n42), .B(n41), .Y(n71) );
  NAND3XLTS U205 ( .A(A[5]), .B(n43), .C(n45), .Y(n44) );
  OAI211XLTS U206 ( .A0(A[5]), .A1(n45), .B0(n71), .C0(n44), .Y(n65) );
  INVX2TS U207 ( .A(n47), .Y(n1553) );
  OAI22X1TS U208 ( .A0(n1554), .A1(n113), .B0(n300), .B1(n1553), .Y(n50) );
  INVX2TS U209 ( .A(B[5]), .Y(n1552) );
  OAI22X1TS U210 ( .A0(n281), .A1(n1552), .B0(n280), .B1(n813), .Y(n49) );
  OAI21XLTS U211 ( .A0(n50), .A1(n49), .B0(n1616), .Y(n48) );
  OAI31X1TS U212 ( .A0(n50), .A1(n1616), .A2(n49), .B0(n48), .Y(n64) );
  INVX2TS U213 ( .A(n53), .Y(Product[5]) );
  OAI22X1TS U214 ( .A0(n1527), .A1(n1660), .B0(n23), .B1(n1659), .Y(n56) );
  INVX2TS U215 ( .A(n15), .Y(n1507) );
  OAI22X1TS U216 ( .A0(n1554), .A1(n1507), .B0(n29), .B1(n1496), .Y(n55) );
  OAI21XLTS U217 ( .A0(n56), .A1(n55), .B0(A[5]), .Y(n54) );
  OAI31X1TS U218 ( .A0(n56), .A1(A[5]), .A2(n55), .B0(n54), .Y(n70) );
  INVX2TS U219 ( .A(A[6]), .Y(n73) );
  OAI22X1TS U220 ( .A0(n14), .A1(A[6]), .B0(n73), .B1(A[5]), .Y(n94) );
  NAND2X1TS U221 ( .A(B[0]), .B(n94), .Y(n76) );
  XOR2XLTS U222 ( .A(n71), .B(n76), .Y(n57) );
  XOR2XLTS U223 ( .A(n70), .B(n57), .Y(n86) );
  INVX2TS U224 ( .A(n59), .Y(n1532) );
  OAI22X1TS U225 ( .A0(n300), .A1(n1532), .B0(n113), .B1(n813), .Y(n62) );
  INVX2TS U226 ( .A(B[6]), .Y(n1533) );
  OAI22X1TS U227 ( .A0(n281), .A1(n1533), .B0(n280), .B1(n1552), .Y(n61) );
  OAI21XLTS U228 ( .A0(n62), .A1(n61), .B0(n1616), .Y(n60) );
  OAI31X1TS U229 ( .A0(n62), .A1(A[2]), .A2(n61), .B0(n60), .Y(n85) );
  INVX2TS U230 ( .A(n66), .Y(Product[6]) );
  OAI22X1TS U231 ( .A0(n29), .A1(n1659), .B0(n1660), .B1(n1537), .Y(n69) );
  OAI22X1TS U232 ( .A0(n1554), .A1(n1496), .B0(n1507), .B1(n813), .Y(n68) );
  OAI21XLTS U233 ( .A0(n69), .A1(n68), .B0(A[5]), .Y(n67) );
  OAI31X1TS U234 ( .A0(n69), .A1(A[5]), .A2(n68), .B0(n67), .Y(n103) );
  AO21XLTS U235 ( .A0(n76), .A1(n71), .B0(n70), .Y(n102) );
  INVX2TS U236 ( .A(n94), .Y(n74) );
  INVX2TS U237 ( .A(A[7]), .Y(n72) );
  OAI22X1TS U238 ( .A0(n1674), .A1(n72), .B0(A[7]), .B1(A[8]), .Y(n95) );
  NOR2XLTS U239 ( .A(n74), .B(n95), .Y(n1333) );
  INVX2TS U240 ( .A(n1333), .Y(n1657) );
  OAI22X1TS U241 ( .A0(n73), .A1(A[7]), .B0(n72), .B1(A[6]), .Y(n93) );
  NAND2X1TS U242 ( .A(n93), .B(n74), .Y(n1322) );
  INVX2TS U243 ( .A(n1322), .Y(n1334) );
  INVX2TS U244 ( .A(n1334), .Y(n1528) );
  OAI222X1TS U245 ( .A0(n1657), .A1(n1516), .B0(n1279), .B1(n23), .C0(n9), 
        .C1(n1528), .Y(n78) );
  INVX2TS U246 ( .A(n78), .Y(n75) );
  NAND3XLTS U247 ( .A(A[8]), .B(n75), .C(n76), .Y(n99) );
  NAND3BXLTS U248 ( .AN(n76), .B(A[8]), .C(n78), .Y(n77) );
  OAI211XLTS U249 ( .A0(A[8]), .A1(n78), .B0(n99), .C0(n77), .Y(n101) );
  INVX2TS U250 ( .A(n80), .Y(n1505) );
  OAI22X1TS U251 ( .A0(n300), .A1(n1505), .B0(n113), .B1(n1552), .Y(n83) );
  INVX2TS U252 ( .A(B[7]), .Y(n1506) );
  OAI22X1TS U253 ( .A0(n281), .A1(n1506), .B0(n280), .B1(n1533), .Y(n82) );
  OAI21XLTS U254 ( .A0(n83), .A1(n82), .B0(n1616), .Y(n81) );
  OAI31X1TS U255 ( .A0(n83), .A1(A[2]), .A2(n82), .B0(n81), .Y(n108) );
  INVX2TS U256 ( .A(n87), .Y(Product[7]) );
  INVX2TS U257 ( .A(n89), .Y(n1500) );
  OAI22X1TS U258 ( .A0(n300), .A1(n1500), .B0(n113), .B1(n1533), .Y(n92) );
  INVX2TS U259 ( .A(B[8]), .Y(n1501) );
  OAI22X1TS U260 ( .A0(n281), .A1(n1501), .B0(n280), .B1(n1506), .Y(n91) );
  OAI21XLTS U261 ( .A0(n92), .A1(n91), .B0(n1616), .Y(n90) );
  OAI31X1TS U262 ( .A0(n92), .A1(A[2]), .A2(n91), .B0(n90), .Y(n124) );
  NOR3XLTS U263 ( .A(n95), .B(n94), .C(n93), .Y(n1332) );
  INVX2TS U264 ( .A(n1332), .Y(n1656) );
  OAI22X1TS U265 ( .A0(n9), .A1(n1656), .B0(n1517), .B1(n1657), .Y(n98) );
  OAI22X1TS U266 ( .A0(n29), .A1(n1279), .B0(n23), .B1(n1528), .Y(n97) );
  OAI21XLTS U267 ( .A0(n98), .A1(n97), .B0(A[8]), .Y(n96) );
  OAI31X1TS U268 ( .A0(n98), .A1(A[8]), .A2(n97), .B0(n96), .Y(n100) );
  NOR2XLTS U269 ( .A(n100), .B(n99), .Y(\mult_x_1/n798 ) );
  AO21XLTS U270 ( .A0(n100), .A1(n99), .B0(\mult_x_1/n798 ), .Y(n1599) );
  OAI22X1TS U271 ( .A0(n1554), .A1(n1659), .B0(n1660), .B1(n1553), .Y(n106) );
  OAI22X1TS U272 ( .A0(n1496), .A1(n813), .B0(n1507), .B1(n1552), .Y(n105) );
  OAI21XLTS U273 ( .A0(n106), .A1(n105), .B0(A[5]), .Y(n104) );
  OAI31X1TS U274 ( .A0(n106), .A1(A[5]), .A2(n105), .B0(n104), .Y(n1597) );
  INVX2TS U275 ( .A(n110), .Y(Product[8]) );
  INVX2TS U276 ( .A(\mult_x_1/n788 ), .Y(n137) );
  INVX2TS U277 ( .A(n112), .Y(n1405) );
  OAI22X1TS U278 ( .A0(n300), .A1(n1405), .B0(n113), .B1(n1501), .Y(n116) );
  INVX2TS U279 ( .A(B[10]), .Y(n1413) );
  INVX2TS U280 ( .A(B[9]), .Y(n1419) );
  OAI22X1TS U281 ( .A0(n281), .A1(n1413), .B0(n280), .B1(n1419), .Y(n115) );
  OAI21XLTS U282 ( .A0(n116), .A1(n115), .B0(n1616), .Y(n114) );
  OAI31X1TS U283 ( .A0(n116), .A1(A[2]), .A2(n115), .B0(n114), .Y(n136) );
  INVX2TS U284 ( .A(\mult_x_1/n793 ), .Y(n128) );
  INVX2TS U285 ( .A(n118), .Y(n1418) );
  OAI22X1TS U286 ( .A0(n300), .A1(n1418), .B0(n113), .B1(n1506), .Y(n121) );
  OAI22X1TS U287 ( .A0(n281), .A1(n1419), .B0(n280), .B1(n1501), .Y(n120) );
  OAI21XLTS U288 ( .A0(n121), .A1(n120), .B0(n1616), .Y(n119) );
  OAI31X1TS U289 ( .A0(n121), .A1(A[2]), .A2(n120), .B0(n119), .Y(n127) );
  INVX2TS U290 ( .A(n125), .Y(Product[10]) );
  INVX2TS U291 ( .A(n129), .Y(Product[9]) );
  INVX2TS U292 ( .A(\mult_x_1/n783 ), .Y(n146) );
  INVX2TS U293 ( .A(n131), .Y(n1409) );
  OAI22X1TS U294 ( .A0(n300), .A1(n1409), .B0(n113), .B1(n1419), .Y(n134) );
  INVX2TS U295 ( .A(B[11]), .Y(n1435) );
  OAI22X1TS U296 ( .A0(n281), .A1(n1435), .B0(n280), .B1(n1413), .Y(n133) );
  OAI21XLTS U297 ( .A0(n134), .A1(n133), .B0(n1616), .Y(n132) );
  OAI31X1TS U298 ( .A0(n134), .A1(A[2]), .A2(n133), .B0(n132), .Y(n145) );
  INVX2TS U299 ( .A(n138), .Y(Product[11]) );
  INVX2TS U300 ( .A(\mult_x_1/n776 ), .Y(n155) );
  INVX2TS U301 ( .A(n140), .Y(n1414) );
  OAI22X1TS U302 ( .A0(n300), .A1(n1414), .B0(n113), .B1(n1413), .Y(n143) );
  INVX2TS U303 ( .A(B[12]), .Y(n1468) );
  OAI22X1TS U304 ( .A0(n281), .A1(n1468), .B0(n280), .B1(n1435), .Y(n142) );
  OAI21XLTS U305 ( .A0(n143), .A1(n142), .B0(n1616), .Y(n141) );
  OAI31X1TS U306 ( .A0(n143), .A1(n1616), .A2(n142), .B0(n141), .Y(n154) );
  INVX2TS U307 ( .A(n147), .Y(Product[12]) );
  INVX2TS U308 ( .A(\mult_x_1/n769 ), .Y(n164) );
  INVX2TS U309 ( .A(n149), .Y(n1436) );
  OAI22X1TS U310 ( .A0(n300), .A1(n1436), .B0(n113), .B1(n1435), .Y(n152) );
  INVX2TS U311 ( .A(B[13]), .Y(n1470) );
  OAI22X1TS U312 ( .A0(n281), .A1(n1470), .B0(n280), .B1(n1468), .Y(n151) );
  OAI21XLTS U313 ( .A0(n152), .A1(n151), .B0(n1616), .Y(n150) );
  OAI31X1TS U314 ( .A0(n152), .A1(A[2]), .A2(n151), .B0(n150), .Y(n163) );
  INVX2TS U315 ( .A(n156), .Y(Product[13]) );
  INVX2TS U316 ( .A(\mult_x_1/n762 ), .Y(n173) );
  INVX2TS U317 ( .A(n158), .Y(n1469) );
  OAI22X1TS U318 ( .A0(n300), .A1(n1469), .B0(n113), .B1(n1468), .Y(n161) );
  INVX2TS U319 ( .A(B[14]), .Y(n1479) );
  OAI22X1TS U320 ( .A0(n281), .A1(n1479), .B0(n280), .B1(n1470), .Y(n160) );
  OAI21XLTS U321 ( .A0(n161), .A1(n160), .B0(n1616), .Y(n159) );
  OAI31X1TS U322 ( .A0(n161), .A1(A[2]), .A2(n160), .B0(n159), .Y(n172) );
  INVX2TS U323 ( .A(n165), .Y(Product[14]) );
  INVX2TS U324 ( .A(\mult_x_1/n754 ), .Y(n182) );
  INVX2TS U325 ( .A(n167), .Y(n1444) );
  OAI22X1TS U326 ( .A0(n300), .A1(n1444), .B0(n113), .B1(n1470), .Y(n170) );
  INVX2TS U327 ( .A(B[15]), .Y(n1482) );
  OAI22X1TS U328 ( .A0(n281), .A1(n1482), .B0(n280), .B1(n1479), .Y(n169) );
  OAI21XLTS U329 ( .A0(n170), .A1(n169), .B0(n1616), .Y(n168) );
  OAI31X1TS U330 ( .A0(n170), .A1(n1616), .A2(n169), .B0(n168), .Y(n181) );
  INVX2TS U331 ( .A(n174), .Y(Product[15]) );
  INVX2TS U332 ( .A(\mult_x_1/n746 ), .Y(n191) );
  INVX2TS U333 ( .A(n176), .Y(n1480) );
  OAI22X1TS U334 ( .A0(n300), .A1(n1480), .B0(n113), .B1(n1479), .Y(n179) );
  INVX2TS U335 ( .A(B[16]), .Y(n1481) );
  OAI22X1TS U336 ( .A0(n281), .A1(n1481), .B0(n280), .B1(n1482), .Y(n178) );
  OAI21XLTS U337 ( .A0(n179), .A1(n178), .B0(n1616), .Y(n177) );
  OAI31X1TS U338 ( .A0(n179), .A1(A[2]), .A2(n178), .B0(n177), .Y(n190) );
  INVX2TS U339 ( .A(n183), .Y(Product[16]) );
  INVX2TS U340 ( .A(\mult_x_1/n738 ), .Y(n200) );
  INVX2TS U341 ( .A(n185), .Y(n1448) );
  OAI22X1TS U342 ( .A0(n300), .A1(n1448), .B0(n113), .B1(n1482), .Y(n188) );
  INVX2TS U343 ( .A(B[17]), .Y(n1449) );
  OAI22X1TS U344 ( .A0(n281), .A1(n1449), .B0(n280), .B1(n1481), .Y(n187) );
  OAI21XLTS U345 ( .A0(n188), .A1(n187), .B0(n1616), .Y(n186) );
  OAI31X1TS U346 ( .A0(n188), .A1(n1616), .A2(n187), .B0(n186), .Y(n199) );
  INVX2TS U347 ( .A(n192), .Y(Product[17]) );
  INVX2TS U348 ( .A(\mult_x_1/n728 ), .Y(n209) );
  INVX2TS U349 ( .A(n194), .Y(n1423) );
  OAI22X1TS U350 ( .A0(n300), .A1(n1423), .B0(n113), .B1(n1481), .Y(n197) );
  INVX2TS U351 ( .A(B[18]), .Y(n1458) );
  OAI22X1TS U352 ( .A0(n281), .A1(n1458), .B0(n280), .B1(n1449), .Y(n196) );
  OAI21XLTS U353 ( .A0(n197), .A1(n196), .B0(n1616), .Y(n195) );
  OAI31X1TS U354 ( .A0(n197), .A1(n1616), .A2(n196), .B0(n195), .Y(n208) );
  INVX2TS U355 ( .A(n201), .Y(Product[18]) );
  INVX2TS U356 ( .A(\mult_x_1/n718 ), .Y(n218) );
  INVX2TS U357 ( .A(n203), .Y(n1393) );
  OAI22X1TS U358 ( .A0(n300), .A1(n1393), .B0(n113), .B1(n1449), .Y(n206) );
  INVX2TS U359 ( .A(B[19]), .Y(n1461) );
  OAI22X1TS U360 ( .A0(n281), .A1(n1461), .B0(n280), .B1(n1458), .Y(n205) );
  OAI21XLTS U361 ( .A0(n206), .A1(n205), .B0(n1616), .Y(n204) );
  OAI31X1TS U362 ( .A0(n206), .A1(n1616), .A2(n205), .B0(n204), .Y(n217) );
  INVX2TS U363 ( .A(n210), .Y(Product[19]) );
  INVX2TS U364 ( .A(\mult_x_1/n708 ), .Y(n227) );
  INVX2TS U365 ( .A(n212), .Y(n1459) );
  OAI22X1TS U366 ( .A0(n300), .A1(n1459), .B0(n113), .B1(n1458), .Y(n215) );
  INVX2TS U367 ( .A(B[20]), .Y(n1460) );
  OAI22X1TS U368 ( .A0(n281), .A1(n1460), .B0(n280), .B1(n1461), .Y(n214) );
  OAI21XLTS U369 ( .A0(n215), .A1(n214), .B0(n1616), .Y(n213) );
  OAI31X1TS U370 ( .A0(n215), .A1(n1616), .A2(n214), .B0(n213), .Y(n226) );
  INVX2TS U371 ( .A(n219), .Y(Product[20]) );
  INVX2TS U372 ( .A(\mult_x_1/n697 ), .Y(n287) );
  INVX2TS U373 ( .A(n221), .Y(n1427) );
  OAI22X1TS U374 ( .A0(n300), .A1(n1427), .B0(n113), .B1(n1461), .Y(n224) );
  INVX2TS U375 ( .A(B[21]), .Y(n1492) );
  OAI22X1TS U376 ( .A0(n281), .A1(n1492), .B0(n280), .B1(n1460), .Y(n223) );
  OAI21XLTS U377 ( .A0(n224), .A1(n223), .B0(n1616), .Y(n222) );
  OAI31X1TS U378 ( .A0(n224), .A1(n1616), .A2(n223), .B0(n222), .Y(n286) );
  INVX2TS U379 ( .A(n228), .Y(Product[21]) );
  INVX2TS U380 ( .A(\mult_x_1/n552 ), .Y(n304) );
  NAND2X1TS U381 ( .A(B[31]), .B(n230), .Y(n1662) );
  OAI21XLTS U382 ( .A0(B[31]), .A1(n230), .B0(n1662), .Y(n1653) );
  INVX2TS U383 ( .A(n1653), .Y(n1606) );
  AOI222XLTS U384 ( .A0(n4), .A1(B[31]), .B0(n2), .B1(n1606), .C0(n231), .C1(
        B[30]), .Y(n232) );
  XOR2XLTS U385 ( .A(n232), .B(n1616), .Y(n303) );
  INVX2TS U386 ( .A(\mult_x_1/n566 ), .Y(n496) );
  INVX2TS U387 ( .A(n234), .Y(n1581) );
  INVX2TS U388 ( .A(B[29]), .Y(n1580) );
  OAI22X1TS U389 ( .A0(n300), .A1(n1581), .B0(n113), .B1(n1580), .Y(n237) );
  INVX2TS U390 ( .A(B[31]), .Y(n1664) );
  INVX2TS U391 ( .A(B[30]), .Y(n1650) );
  OAI22X1TS U392 ( .A0(n281), .A1(n1664), .B0(n280), .B1(n1650), .Y(n236) );
  OAI21XLTS U393 ( .A0(n237), .A1(n236), .B0(n1616), .Y(n235) );
  OAI31X1TS U394 ( .A0(n237), .A1(n1616), .A2(n236), .B0(n235), .Y(n495) );
  INVX2TS U395 ( .A(\mult_x_1/n580 ), .Y(n458) );
  INVX2TS U396 ( .A(n239), .Y(n1561) );
  INVX2TS U397 ( .A(B[28]), .Y(n1560) );
  OAI22X1TS U398 ( .A0(n300), .A1(n1561), .B0(n113), .B1(n1560), .Y(n242) );
  OAI22X1TS U399 ( .A0(n281), .A1(n1650), .B0(n280), .B1(n1580), .Y(n241) );
  OAI21XLTS U400 ( .A0(n242), .A1(n241), .B0(n1616), .Y(n240) );
  OAI31X1TS U401 ( .A0(n242), .A1(n1616), .A2(n241), .B0(n240), .Y(n457) );
  INVX2TS U402 ( .A(\mult_x_1/n594 ), .Y(n448) );
  INVX2TS U403 ( .A(n244), .Y(n1440) );
  INVX2TS U404 ( .A(B[27]), .Y(n1454) );
  OAI22X1TS U405 ( .A0(n300), .A1(n1440), .B0(n113), .B1(n1454), .Y(n247) );
  OAI22X1TS U406 ( .A0(n281), .A1(n1580), .B0(n280), .B1(n1560), .Y(n246) );
  OAI21XLTS U407 ( .A0(n247), .A1(n246), .B0(n1616), .Y(n245) );
  OAI31X1TS U408 ( .A0(n247), .A1(A[2]), .A2(n246), .B0(n245), .Y(n447) );
  INVX2TS U409 ( .A(\mult_x_1/n608 ), .Y(n441) );
  INVX2TS U410 ( .A(n249), .Y(n1453) );
  INVX2TS U411 ( .A(B[26]), .Y(n1475) );
  OAI22X1TS U412 ( .A0(n300), .A1(n1453), .B0(n113), .B1(n1475), .Y(n252) );
  OAI22X1TS U413 ( .A0(n281), .A1(n1560), .B0(n280), .B1(n1454), .Y(n251) );
  OAI21XLTS U414 ( .A0(n252), .A1(n251), .B0(n1616), .Y(n250) );
  OAI31X1TS U415 ( .A0(n252), .A1(A[2]), .A2(n251), .B0(n250), .Y(n440) );
  INVX2TS U416 ( .A(\mult_x_1/n622 ), .Y(n369) );
  INVX2TS U417 ( .A(n254), .Y(n1397) );
  INVX2TS U418 ( .A(B[25]), .Y(n1487) );
  OAI22X1TS U419 ( .A0(n300), .A1(n1397), .B0(n113), .B1(n1487), .Y(n257) );
  OAI22X1TS U420 ( .A0(n281), .A1(n1454), .B0(n280), .B1(n1475), .Y(n256) );
  OAI21XLTS U421 ( .A0(n257), .A1(n256), .B0(n1616), .Y(n255) );
  OAI31X1TS U422 ( .A0(n257), .A1(n1616), .A2(n256), .B0(n255), .Y(n368) );
  INVX2TS U423 ( .A(\mult_x_1/n636 ), .Y(n352) );
  INVX2TS U424 ( .A(n259), .Y(n1474) );
  INVX2TS U425 ( .A(B[24]), .Y(n1488) );
  OAI22X1TS U426 ( .A0(n300), .A1(n1474), .B0(n113), .B1(n1488), .Y(n262) );
  OAI22X1TS U427 ( .A0(n281), .A1(n1475), .B0(n280), .B1(n1487), .Y(n261) );
  OAI21XLTS U428 ( .A0(n262), .A1(n261), .B0(n1616), .Y(n260) );
  OAI31X1TS U429 ( .A0(n262), .A1(A[2]), .A2(n261), .B0(n260), .Y(n351) );
  INVX2TS U430 ( .A(\mult_x_1/n649 ), .Y(n365) );
  INVX2TS U431 ( .A(n264), .Y(n1486) );
  INVX2TS U432 ( .A(B[23]), .Y(n1494) );
  OAI22X1TS U433 ( .A0(n300), .A1(n1486), .B0(n113), .B1(n1494), .Y(n267) );
  OAI22X1TS U434 ( .A0(n281), .A1(n1487), .B0(n280), .B1(n1488), .Y(n266) );
  OAI21XLTS U435 ( .A0(n267), .A1(n266), .B0(n1616), .Y(n265) );
  OAI31X1TS U436 ( .A0(n267), .A1(n1616), .A2(n266), .B0(n265), .Y(n364) );
  INVX2TS U437 ( .A(\mult_x_1/n662 ), .Y(n336) );
  INVX2TS U438 ( .A(n269), .Y(n1431) );
  INVX2TS U439 ( .A(B[22]), .Y(n1495) );
  OAI22X1TS U440 ( .A0(n300), .A1(n1431), .B0(n113), .B1(n1495), .Y(n272) );
  OAI22X1TS U441 ( .A0(n281), .A1(n1488), .B0(n280), .B1(n1494), .Y(n271) );
  OAI21XLTS U442 ( .A0(n272), .A1(n271), .B0(n1616), .Y(n270) );
  OAI31X1TS U443 ( .A0(n272), .A1(n1616), .A2(n271), .B0(n270), .Y(n335) );
  INVX2TS U444 ( .A(\mult_x_1/n675 ), .Y(n316) );
  INVX2TS U445 ( .A(n274), .Y(n1493) );
  OAI22X1TS U446 ( .A0(n300), .A1(n1493), .B0(n113), .B1(n1492), .Y(n277) );
  OAI22X1TS U447 ( .A0(n281), .A1(n1494), .B0(n280), .B1(n1495), .Y(n276) );
  OAI21XLTS U448 ( .A0(n277), .A1(n276), .B0(n1616), .Y(n275) );
  OAI31X1TS U449 ( .A0(n277), .A1(n1616), .A2(n276), .B0(n275), .Y(n315) );
  INVX2TS U450 ( .A(\mult_x_1/n686 ), .Y(n308) );
  INVX2TS U451 ( .A(n279), .Y(n1401) );
  OAI22X1TS U452 ( .A0(n300), .A1(n1401), .B0(n113), .B1(n1460), .Y(n284) );
  OAI22X1TS U453 ( .A0(n281), .A1(n1495), .B0(n280), .B1(n1492), .Y(n283) );
  OAI21XLTS U454 ( .A0(n284), .A1(n283), .B0(n1616), .Y(n282) );
  OAI31X1TS U455 ( .A0(n284), .A1(A[2]), .A2(n283), .B0(n282), .Y(n307) );
  INVX2TS U456 ( .A(n288), .Y(Product[32]) );
  INVX2TS U457 ( .A(A[30]), .Y(n290) );
  INVX2TS U458 ( .A(A[29]), .Y(n1625) );
  AOI22X1TS U459 ( .A0(A[29]), .A1(A[30]), .B0(n290), .B1(n1625), .Y(n795) );
  INVX2TS U460 ( .A(A[31]), .Y(n289) );
  NAND2X1TS U461 ( .A(n795), .B(n289), .Y(n1579) );
  AOI221XLTS U462 ( .A0(A[30]), .A1(A[31]), .B0(n290), .B1(n289), .C0(n795), 
        .Y(n291) );
  INVX2TS U463 ( .A(n291), .Y(n1591) );
  NAND2X1TS U464 ( .A(n795), .B(A[31]), .Y(n1663) );
  OAI22X1TS U465 ( .A0(n1453), .A1(n1663), .B0(n1475), .B1(n1559), .Y(n292) );
  AOI21X1TS U466 ( .A0(B[27]), .A1(n1584), .B0(n292), .Y(n293) );
  OAI21XLTS U467 ( .A0(n1560), .A1(n1579), .B0(n293), .Y(\mult_x_1/n916 ) );
  OAI22X1TS U468 ( .A0(n1397), .A1(n1663), .B0(n1487), .B1(n1559), .Y(n294) );
  AOI21X1TS U469 ( .A0(B[26]), .A1(n1584), .B0(n294), .Y(n295) );
  OAI21XLTS U470 ( .A0(n1454), .A1(n1579), .B0(n295), .Y(\mult_x_1/n917 ) );
  OAI22X1TS U471 ( .A0(n1474), .A1(n1663), .B0(n1488), .B1(n1559), .Y(n296) );
  AOI21X1TS U472 ( .A0(B[25]), .A1(n1584), .B0(n296), .Y(n297) );
  OAI21XLTS U473 ( .A0(n1475), .A1(n1579), .B0(n297), .Y(\mult_x_1/n918 ) );
  CLKBUFX2TS U474 ( .A(n1663), .Y(n1592) );
  OAI22X1TS U475 ( .A0(n1486), .A1(n1592), .B0(n1494), .B1(n1559), .Y(n298) );
  AOI21X1TS U476 ( .A0(B[24]), .A1(n1584), .B0(n298), .Y(n299) );
  OAI21XLTS U477 ( .A0(n1487), .A1(n1579), .B0(n299), .Y(n1620) );
  INVX2TS U478 ( .A(\mult_x_1/n307 ), .Y(\mult_x_1/n312 ) );
  INVX2TS U479 ( .A(\mult_x_1/n538 ), .Y(n312) );
  OAI22X1TS U480 ( .A0(n300), .A1(n1662), .B0(n113), .B1(n1664), .Y(n301) );
  XOR2XLTS U481 ( .A(n693), .B(n301), .Y(n311) );
  INVX2TS U482 ( .A(n305), .Y(Product[33]) );
  INVX2TS U483 ( .A(n309), .Y(Product[22]) );
  INVX2TS U484 ( .A(\mult_x_1/n537 ), .Y(n332) );
  INVX2TS U485 ( .A(\mult_x_1/n524 ), .Y(n331) );
  INVX2TS U486 ( .A(n313), .Y(Product[34]) );
  INVX2TS U487 ( .A(n317), .Y(Product[23]) );
  OAI2BB2XLTS U488 ( .B0(n1671), .B1(A[27]), .A0N(A[27]), .A1N(n1671), .Y(n321) );
  INVX2TS U489 ( .A(n321), .Y(n790) );
  OAI2BB2XLTS U490 ( .B0(A[28]), .B1(A[29]), .A0N(A[29]), .A1N(A[28]), .Y(n320) );
  NOR2XLTS U491 ( .A(n790), .B(n320), .Y(n1387) );
  INVX2TS U492 ( .A(n1387), .Y(n1565) );
  XOR2XLTS U493 ( .A(A[27]), .B(A[28]), .Y(n318) );
  NOR3XLTS U494 ( .A(n320), .B(n321), .C(n318), .Y(n1385) );
  INVX2TS U495 ( .A(n1385), .Y(n1564) );
  OAI22X1TS U496 ( .A0(n1565), .A1(n1581), .B0(n1564), .B1(n1580), .Y(n325) );
  NAND2X1TS U497 ( .A(n318), .B(n790), .Y(n319) );
  INVX2TS U498 ( .A(n319), .Y(n1386) );
  OAI22X1TS U499 ( .A0(n319), .A1(n1650), .B0(n322), .B1(n1664), .Y(n324) );
  OAI21XLTS U500 ( .A0(n325), .A1(n324), .B0(n1625), .Y(n323) );
  OAI31X1TS U501 ( .A0(n325), .A1(n1625), .A2(n324), .B0(n323), .Y(
        \mult_x_1/n945 ) );
  OAI22X1TS U502 ( .A0(n1401), .A1(n1592), .B0(n1460), .B1(n1559), .Y(n326) );
  AOI21X1TS U503 ( .A0(B[21]), .A1(n1584), .B0(n326), .Y(n327) );
  OAI21XLTS U504 ( .A0(n1495), .A1(n1579), .B0(n327), .Y(\mult_x_1/n922 ) );
  OAI22X1TS U505 ( .A0(n1427), .A1(n1592), .B0(n1461), .B1(n1559), .Y(n328) );
  AOI21X1TS U506 ( .A0(B[20]), .A1(n1584), .B0(n328), .Y(n329) );
  OAI21XLTS U507 ( .A0(n1492), .A1(n1579), .B0(n329), .Y(\mult_x_1/n923 ) );
  INVX2TS U508 ( .A(\mult_x_1/n523 ), .Y(n361) );
  INVX2TS U509 ( .A(\mult_x_1/n510 ), .Y(n360) );
  INVX2TS U510 ( .A(n333), .Y(Product[35]) );
  INVX2TS U511 ( .A(n337), .Y(Product[24]) );
  OAI22X1TS U512 ( .A0(n1565), .A1(n1440), .B0(n1564), .B1(n1454), .Y(n340) );
  OAI22X1TS U513 ( .A0(n796), .A1(n1560), .B0(n322), .B1(n1580), .Y(n339) );
  OAI21XLTS U514 ( .A0(n340), .A1(n339), .B0(n1625), .Y(n338) );
  OAI31X1TS U515 ( .A0(n340), .A1(n1625), .A2(n339), .B0(n338), .Y(
        \mult_x_1/n947 ) );
  OAI22X1TS U516 ( .A0(n1565), .A1(n1561), .B0(n1564), .B1(n1560), .Y(n343) );
  OAI22X1TS U517 ( .A0(n319), .A1(n1580), .B0(n322), .B1(n1650), .Y(n342) );
  OAI21XLTS U518 ( .A0(n343), .A1(n342), .B0(n1625), .Y(n341) );
  OAI31X1TS U519 ( .A0(n343), .A1(n1625), .A2(n342), .B0(n341), .Y(
        \mult_x_1/n946 ) );
  INVX2TS U520 ( .A(\mult_x_1/n366 ), .Y(n372) );
  NOR2XLTS U521 ( .A(n1461), .B(n1579), .Y(n345) );
  OAI22X1TS U522 ( .A0(n1393), .A1(n1592), .B0(n1449), .B1(n1559), .Y(n344) );
  AOI211XLTS U523 ( .A0(n1584), .A1(B[18]), .B0(n345), .C0(n344), .Y(n371) );
  INVX2TS U524 ( .A(n346), .Y(\mult_x_1/n356 ) );
  OAI22X1TS U525 ( .A0(n1565), .A1(n1453), .B0(n1564), .B1(n1475), .Y(n349) );
  OAI22X1TS U526 ( .A0(n796), .A1(n1454), .B0(n322), .B1(n1560), .Y(n348) );
  OAI21XLTS U527 ( .A0(n349), .A1(n348), .B0(n1625), .Y(n347) );
  OAI31X1TS U528 ( .A0(n349), .A1(n1625), .A2(n348), .B0(n347), .Y(
        \mult_x_1/n948 ) );
  INVX2TS U529 ( .A(n353), .Y(Product[26]) );
  OAI22X1TS U530 ( .A0(n1459), .A1(n1592), .B0(n1458), .B1(n1559), .Y(n354) );
  AOI21X1TS U531 ( .A0(B[19]), .A1(n1584), .B0(n354), .Y(n355) );
  OAI21XLTS U532 ( .A0(n1460), .A1(n1579), .B0(n355), .Y(\mult_x_1/n341 ) );
  INVX2TS U533 ( .A(\mult_x_1/n341 ), .Y(\mult_x_1/n349 ) );
  OAI22X1TS U534 ( .A0(n1565), .A1(n1397), .B0(n1564), .B1(n1487), .Y(n358) );
  OAI22X1TS U535 ( .A0(n796), .A1(n1475), .B0(n322), .B1(n1454), .Y(n357) );
  OAI21XLTS U536 ( .A0(n358), .A1(n357), .B0(n1625), .Y(n356) );
  OAI31X1TS U537 ( .A0(n358), .A1(n1625), .A2(n357), .B0(n356), .Y(
        \mult_x_1/n949 ) );
  INVX2TS U538 ( .A(\mult_x_1/n509 ), .Y(n387) );
  INVX2TS U539 ( .A(\mult_x_1/n496 ), .Y(n386) );
  INVX2TS U540 ( .A(n362), .Y(Product[36]) );
  INVX2TS U541 ( .A(n366), .Y(Product[25]) );
  INVX2TS U542 ( .A(n370), .Y(Product[27]) );
  INVX2TS U543 ( .A(n373), .Y(\mult_x_1/n357 ) );
  OAI22X1TS U544 ( .A0(n1565), .A1(n1474), .B0(n1564), .B1(n1488), .Y(n376) );
  OAI22X1TS U545 ( .A0(n796), .A1(n1487), .B0(n322), .B1(n1475), .Y(n375) );
  OAI21XLTS U546 ( .A0(n376), .A1(n375), .B0(A[29]), .Y(n374) );
  OAI31X1TS U547 ( .A0(n376), .A1(A[29]), .A2(n375), .B0(n374), .Y(n399) );
  NOR2XLTS U548 ( .A(n1494), .B(n1579), .Y(n378) );
  OAI22X1TS U549 ( .A0(n1493), .A1(n1592), .B0(n1492), .B1(n1559), .Y(n377) );
  AOI211XLTS U550 ( .A0(n1584), .A1(B[22]), .B0(n378), .C0(n377), .Y(n398) );
  NOR2XLTS U551 ( .A(n1488), .B(n1579), .Y(n380) );
  OAI22X1TS U552 ( .A0(n1431), .A1(n1592), .B0(n1495), .B1(n1559), .Y(n379) );
  AOI211XLTS U553 ( .A0(B[23]), .A1(n1584), .B0(n380), .C0(n379), .Y(n418) );
  INVX2TS U554 ( .A(n381), .Y(\mult_x_1/n320 ) );
  OAI22X1TS U555 ( .A0(n1565), .A1(n1486), .B0(n1564), .B1(n1494), .Y(n384) );
  OAI22X1TS U556 ( .A0(n796), .A1(n1488), .B0(n322), .B1(n1487), .Y(n383) );
  OAI21XLTS U557 ( .A0(n384), .A1(n383), .B0(n1625), .Y(n382) );
  OAI31X1TS U558 ( .A0(n384), .A1(n1625), .A2(n383), .B0(n382), .Y(
        \mult_x_1/n951 ) );
  INVX2TS U559 ( .A(\mult_x_1/n495 ), .Y(n407) );
  INVX2TS U560 ( .A(\mult_x_1/n482 ), .Y(n406) );
  INVX2TS U561 ( .A(n388), .Y(Product[37]) );
  INVX2TS U562 ( .A(A[24]), .Y(n389) );
  OAI22X1TS U563 ( .A0(n1621), .A1(A[24]), .B0(n389), .B1(A[23]), .Y(n393) );
  INVX2TS U564 ( .A(n393), .Y(n895) );
  INVX2TS U565 ( .A(A[25]), .Y(n390) );
  OAI22X1TS U566 ( .A0(n1671), .A1(n390), .B0(A[25]), .B1(A[26]), .Y(n392) );
  NOR2XLTS U567 ( .A(n895), .B(n392), .Y(n434) );
  INVX2TS U568 ( .A(n434), .Y(n1602) );
  AOI22X1TS U569 ( .A0(A[24]), .A1(A[25]), .B0(n390), .B1(n389), .Y(n391) );
  NOR3XLTS U570 ( .A(n392), .B(n393), .C(n391), .Y(n432) );
  INVX2TS U571 ( .A(n432), .Y(n1601) );
  OAI22X1TS U572 ( .A0(n1602), .A1(n1581), .B0(n1601), .B1(n1580), .Y(n397) );
  NAND2X1TS U573 ( .A(n391), .B(n895), .Y(n896) );
  INVX2TS U574 ( .A(n896), .Y(n433) );
  INVX2TS U575 ( .A(n433), .Y(n927) );
  NAND2X1TS U576 ( .A(n393), .B(n392), .Y(n394) );
  INVX2TS U577 ( .A(n394), .Y(n899) );
  OAI22X1TS U578 ( .A0(n927), .A1(n1650), .B0(n902), .B1(n1664), .Y(n396) );
  OAI21XLTS U579 ( .A0(n397), .A1(n396), .B0(n1671), .Y(n395) );
  OAI31X1TS U580 ( .A0(n397), .A1(n1671), .A2(n396), .B0(n395), .Y(
        \mult_x_1/n980 ) );
  INVX2TS U581 ( .A(n400), .Y(\mult_x_1/n328 ) );
  OAI22X1TS U582 ( .A0(n1480), .A1(n1592), .B0(n1479), .B1(n1559), .Y(n401) );
  AOI21X1TS U583 ( .A0(B[15]), .A1(n1584), .B0(n401), .Y(n402) );
  OAI21XLTS U584 ( .A0(n1481), .A1(n1579), .B0(n402), .Y(\mult_x_1/n927 ) );
  OAI22X1TS U585 ( .A0(n1444), .A1(n1592), .B0(n1470), .B1(n1559), .Y(n403) );
  AOI21X1TS U586 ( .A0(B[14]), .A1(n1584), .B0(n403), .Y(n404) );
  OAI21XLTS U587 ( .A0(n1482), .A1(n1579), .B0(n404), .Y(\mult_x_1/n928 ) );
  INVX2TS U588 ( .A(\mult_x_1/n481 ), .Y(n468) );
  INVX2TS U589 ( .A(\mult_x_1/n469 ), .Y(n467) );
  INVX2TS U590 ( .A(n408), .Y(Product[38]) );
  OAI22X1TS U591 ( .A0(n1565), .A1(n1431), .B0(n1564), .B1(n1495), .Y(n411) );
  OAI22X1TS U592 ( .A0(n796), .A1(n1494), .B0(n322), .B1(n1488), .Y(n410) );
  OAI21XLTS U593 ( .A0(n411), .A1(n410), .B0(n1625), .Y(n409) );
  OAI31X1TS U594 ( .A0(n411), .A1(n1625), .A2(n410), .B0(n409), .Y(
        \mult_x_1/n952 ) );
  OAI22X1TS U595 ( .A0(n1565), .A1(n1493), .B0(n1564), .B1(n1492), .Y(n414) );
  OAI22X1TS U596 ( .A0(n796), .A1(n1495), .B0(n322), .B1(n1494), .Y(n413) );
  OAI21XLTS U597 ( .A0(n414), .A1(n413), .B0(n1625), .Y(n412) );
  OAI31X1TS U598 ( .A0(n414), .A1(n1625), .A2(n413), .B0(n412), .Y(
        \mult_x_1/n953 ) );
  INVX2TS U599 ( .A(\mult_x_1/n428 ), .Y(n471) );
  INVX2TS U600 ( .A(n1591), .Y(n1584) );
  NOR2XLTS U601 ( .A(n1470), .B(n1579), .Y(n416) );
  OAI22X1TS U602 ( .A0(n1436), .A1(n1592), .B0(n1435), .B1(n1559), .Y(n415) );
  AOI211XLTS U603 ( .A0(n1584), .A1(B[12]), .B0(n416), .C0(n415), .Y(n470) );
  INVX2TS U604 ( .A(n417), .Y(\mult_x_1/n415 ) );
  INVX2TS U605 ( .A(n420), .Y(\mult_x_1/n321 ) );
  OAI22X1TS U606 ( .A0(n1565), .A1(n1401), .B0(n1564), .B1(n1460), .Y(n423) );
  OAI22X1TS U607 ( .A0(n319), .A1(n1492), .B0(n322), .B1(n1495), .Y(n422) );
  OAI21XLTS U608 ( .A0(n423), .A1(n422), .B0(n1625), .Y(n421) );
  OAI31X1TS U609 ( .A0(n423), .A1(n1625), .A2(n422), .B0(n421), .Y(
        \mult_x_1/n954 ) );
  OAI22X1TS U610 ( .A0(n1602), .A1(n1561), .B0(n1601), .B1(n1560), .Y(n426) );
  OAI22X1TS U611 ( .A0(n927), .A1(n1580), .B0(n902), .B1(n1650), .Y(n425) );
  OAI21XLTS U612 ( .A0(n426), .A1(n425), .B0(n1671), .Y(n424) );
  OAI31X1TS U613 ( .A0(n426), .A1(n1671), .A2(n425), .B0(n424), .Y(
        \mult_x_1/n981 ) );
  OAI22X1TS U614 ( .A0(n1602), .A1(n1440), .B0(n1601), .B1(n1454), .Y(n429) );
  OAI22X1TS U615 ( .A0(n927), .A1(n1560), .B0(n902), .B1(n1580), .Y(n428) );
  OAI21XLTS U616 ( .A0(n429), .A1(n428), .B0(n1671), .Y(n427) );
  OAI31X1TS U617 ( .A0(n429), .A1(n1671), .A2(n428), .B0(n427), .Y(
        \mult_x_1/n982 ) );
  OAI22X1TS U618 ( .A0(n1469), .A1(n1592), .B0(n1468), .B1(n1559), .Y(n430) );
  AOI21X1TS U619 ( .A0(B[13]), .A1(n1584), .B0(n430), .Y(n431) );
  OAI21XLTS U620 ( .A0(n1479), .A1(n1579), .B0(n431), .Y(\mult_x_1/n394 ) );
  INVX2TS U621 ( .A(\mult_x_1/n394 ), .Y(\mult_x_1/n405 ) );
  AOI222XLTS U622 ( .A0(n434), .A1(n1606), .B0(n433), .B1(B[31]), .C0(n432), 
        .C1(B[30]), .Y(n435) );
  XOR2XLTS U623 ( .A(n1671), .B(n435), .Y(\mult_x_1/n979 ) );
  OAI22X1TS U624 ( .A0(n1602), .A1(n1453), .B0(n1601), .B1(n1475), .Y(n438) );
  OAI22X1TS U625 ( .A0(n927), .A1(n1454), .B0(n902), .B1(n1560), .Y(n437) );
  OAI21XLTS U626 ( .A0(n438), .A1(n437), .B0(n1671), .Y(n436) );
  OAI31X1TS U627 ( .A0(n438), .A1(n1671), .A2(n437), .B0(n436), .Y(
        \mult_x_1/n983 ) );
  INVX2TS U628 ( .A(n442), .Y(Product[28]) );
  OAI22X1TS U629 ( .A0(n1602), .A1(n1397), .B0(n1601), .B1(n1487), .Y(n445) );
  OAI22X1TS U630 ( .A0(n927), .A1(n1475), .B0(n394), .B1(n1454), .Y(n444) );
  OAI21XLTS U631 ( .A0(n445), .A1(n444), .B0(n1671), .Y(n443) );
  OAI31X1TS U632 ( .A0(n445), .A1(n1671), .A2(n444), .B0(n443), .Y(
        \mult_x_1/n984 ) );
  INVX2TS U633 ( .A(n449), .Y(Product[29]) );
  OAI22X1TS U634 ( .A0(n1565), .A1(n1427), .B0(n1564), .B1(n1461), .Y(n452) );
  INVX2TS U635 ( .A(n1386), .Y(n796) );
  OAI22X1TS U636 ( .A0(n796), .A1(n1460), .B0(n322), .B1(n1492), .Y(n451) );
  OAI21XLTS U637 ( .A0(n452), .A1(n451), .B0(A[29]), .Y(n450) );
  OAI31X1TS U638 ( .A0(n452), .A1(A[29]), .A2(n451), .B0(n450), .Y(n490) );
  NOR2XLTS U639 ( .A(n1458), .B(n1579), .Y(n454) );
  OAI22X1TS U640 ( .A0(n1423), .A1(n1592), .B0(n1481), .B1(n1559), .Y(n453) );
  AOI211XLTS U641 ( .A0(n1584), .A1(B[17]), .B0(n454), .C0(n453), .Y(n489) );
  INVX2TS U642 ( .A(n455), .Y(\mult_x_1/n364 ) );
  INVX2TS U643 ( .A(n459), .Y(Product[30]) );
  OAI22X1TS U644 ( .A0(n1565), .A1(n1459), .B0(n1564), .B1(n1458), .Y(n462) );
  OAI22X1TS U645 ( .A0(n796), .A1(n1461), .B0(n322), .B1(n1460), .Y(n461) );
  OAI21XLTS U646 ( .A0(n462), .A1(n461), .B0(A[29]), .Y(n460) );
  OAI31X1TS U647 ( .A0(n462), .A1(A[29]), .A2(n461), .B0(n460), .Y(n487) );
  NOR2XLTS U648 ( .A(n1449), .B(n1579), .Y(n464) );
  OAI22X1TS U649 ( .A0(n1448), .A1(n1592), .B0(n1482), .B1(n1559), .Y(n463) );
  AOI211XLTS U650 ( .A0(n1584), .A1(B[16]), .B0(n464), .C0(n463), .Y(n486) );
  INVX2TS U651 ( .A(n465), .Y(\mult_x_1/n374 ) );
  INVX2TS U652 ( .A(\mult_x_1/n468 ), .Y(n484) );
  INVX2TS U653 ( .A(\mult_x_1/n455 ), .Y(n483) );
  INVX2TS U654 ( .A(n469), .Y(Product[39]) );
  INVX2TS U655 ( .A(n472), .Y(\mult_x_1/n416 ) );
  OAI22X1TS U656 ( .A0(n1565), .A1(n1393), .B0(n1564), .B1(n1449), .Y(n475) );
  OAI22X1TS U657 ( .A0(n319), .A1(n1458), .B0(n322), .B1(n1461), .Y(n474) );
  OAI21XLTS U658 ( .A0(n475), .A1(n474), .B0(n1625), .Y(n473) );
  OAI31X1TS U659 ( .A0(n475), .A1(n1625), .A2(n474), .B0(n473), .Y(
        \mult_x_1/n957 ) );
  OAI22X1TS U660 ( .A0(n1602), .A1(n1474), .B0(n1601), .B1(n1488), .Y(n478) );
  OAI22X1TS U661 ( .A0(n927), .A1(n1487), .B0(n394), .B1(n1475), .Y(n477) );
  OAI21XLTS U662 ( .A0(n478), .A1(n477), .B0(n1671), .Y(n476) );
  OAI31X1TS U663 ( .A0(n478), .A1(n1671), .A2(n477), .B0(n476), .Y(
        \mult_x_1/n985 ) );
  OAI22X1TS U664 ( .A0(n1602), .A1(n1486), .B0(n1601), .B1(n1494), .Y(n481) );
  OAI22X1TS U665 ( .A0(n927), .A1(n1488), .B0(n394), .B1(n1487), .Y(n480) );
  OAI21XLTS U666 ( .A0(n481), .A1(n480), .B0(n1671), .Y(n479) );
  OAI31X1TS U667 ( .A0(n481), .A1(n1671), .A2(n480), .B0(n479), .Y(
        \mult_x_1/n986 ) );
  INVX2TS U668 ( .A(\mult_x_1/n454 ), .Y(n517) );
  INVX2TS U669 ( .A(\mult_x_1/n444 ), .Y(n516) );
  INVX2TS U670 ( .A(n485), .Y(Product[40]) );
  INVX2TS U671 ( .A(n488), .Y(\mult_x_1/n375 ) );
  INVX2TS U672 ( .A(n491), .Y(\mult_x_1/n365 ) );
  OAI22X1TS U673 ( .A0(n1418), .A1(n1592), .B0(n1506), .B1(n1559), .Y(n492) );
  AOI21X1TS U674 ( .A0(B[8]), .A1(n1584), .B0(n492), .Y(n493) );
  OAI21XLTS U675 ( .A0(n1419), .A1(n1579), .B0(n493), .Y(\mult_x_1/n933 ) );
  INVX2TS U676 ( .A(n497), .Y(Product[31]) );
  AOI2BB2XLTS U677 ( .B0(A[23]), .B1(A[22]), .A0N(A[22]), .A1N(A[23]), .Y(n500) );
  OAI2BB2XLTS U678 ( .B0(n1672), .B1(A[21]), .A0N(A[21]), .A1N(n1672), .Y(n498) );
  OAI22X1TS U679 ( .A0(n723), .A1(n1581), .B0(n727), .B1(n1664), .Y(n503) );
  XNOR2X1TS U680 ( .A(A[22]), .B(A[21]), .Y(n499) );
  INVX2TS U681 ( .A(n498), .Y(n1012) );
  NAND3XLTS U682 ( .A(n500), .B(n1012), .C(n499), .Y(n1642) );
  CLKBUFX2TS U683 ( .A(n1642), .Y(n1640) );
  OAI22X1TS U684 ( .A0(n1643), .A1(n1650), .B0(n1640), .B1(n1580), .Y(n502) );
  OAI21XLTS U685 ( .A0(n503), .A1(n502), .B0(n1621), .Y(n501) );
  OAI31X1TS U686 ( .A0(n503), .A1(n1621), .A2(n502), .B0(n501), .Y(
        \mult_x_1/n1015 ) );
  OAI22X1TS U687 ( .A0(n1405), .A1(n1592), .B0(n1501), .B1(n1559), .Y(n504) );
  AOI21X1TS U688 ( .A0(B[9]), .A1(n1584), .B0(n504), .Y(n505) );
  OAI21XLTS U689 ( .A0(n1413), .A1(n1579), .B0(n505), .Y(\mult_x_1/n932 ) );
  OAI22X1TS U690 ( .A0(n1565), .A1(n1448), .B0(n1564), .B1(n1482), .Y(n508) );
  OAI22X1TS U691 ( .A0(n319), .A1(n1481), .B0(n322), .B1(n1449), .Y(n507) );
  OAI21XLTS U692 ( .A0(n508), .A1(n507), .B0(n1625), .Y(n506) );
  OAI31X1TS U693 ( .A0(n508), .A1(n1625), .A2(n507), .B0(n506), .Y(
        \mult_x_1/n959 ) );
  OAI22X1TS U694 ( .A0(n1565), .A1(n1423), .B0(n1564), .B1(n1481), .Y(n511) );
  OAI22X1TS U695 ( .A0(n319), .A1(n1449), .B0(n322), .B1(n1458), .Y(n510) );
  OAI21XLTS U696 ( .A0(n511), .A1(n510), .B0(n1625), .Y(n509) );
  OAI31X1TS U697 ( .A0(n511), .A1(n1625), .A2(n510), .B0(n509), .Y(
        \mult_x_1/n958 ) );
  NOR2XLTS U698 ( .A(n1506), .B(n1579), .Y(n513) );
  OAI22X1TS U699 ( .A0(n1505), .A1(n1592), .B0(n1552), .B1(n1559), .Y(n512) );
  AOI211XLTS U700 ( .A0(n1584), .A1(B[6]), .B0(n513), .C0(n512), .Y(n571) );
  INVX2TS U701 ( .A(n514), .Y(\mult_x_1/n492 ) );
  INVX2TS U702 ( .A(\mult_x_1/n443 ), .Y(n569) );
  INVX2TS U703 ( .A(\mult_x_1/n432 ), .Y(n568) );
  INVX2TS U704 ( .A(n518), .Y(Product[41]) );
  OAI22X1TS U705 ( .A0(n1500), .A1(n1592), .B0(n1533), .B1(n1559), .Y(n519) );
  AOI21X1TS U706 ( .A0(B[7]), .A1(n1584), .B0(n519), .Y(n520) );
  OAI21XLTS U707 ( .A0(n1501), .A1(n1579), .B0(n520), .Y(\mult_x_1/n465 ) );
  INVX2TS U708 ( .A(\mult_x_1/n465 ), .Y(\mult_x_1/n479 ) );
  OAI22X1TS U709 ( .A0(n1602), .A1(n1431), .B0(n1601), .B1(n1495), .Y(n523) );
  OAI22X1TS U710 ( .A0(n927), .A1(n1494), .B0(n394), .B1(n1488), .Y(n522) );
  OAI21XLTS U711 ( .A0(n523), .A1(n522), .B0(n1671), .Y(n521) );
  OAI31X1TS U712 ( .A0(n523), .A1(n1671), .A2(n522), .B0(n521), .Y(
        \mult_x_1/n987 ) );
  OAI22X1TS U713 ( .A0(n1602), .A1(n1493), .B0(n1601), .B1(n1492), .Y(n526) );
  OAI22X1TS U714 ( .A0(n927), .A1(n1495), .B0(n394), .B1(n1494), .Y(n525) );
  OAI21XLTS U715 ( .A0(n526), .A1(n525), .B0(n1671), .Y(n524) );
  OAI31X1TS U716 ( .A0(n526), .A1(n1671), .A2(n525), .B0(n524), .Y(
        \mult_x_1/n988 ) );
  OAI22X1TS U717 ( .A0(n1565), .A1(n1480), .B0(n1564), .B1(n1479), .Y(n529) );
  OAI22X1TS U718 ( .A0(n319), .A1(n1482), .B0(n322), .B1(n1481), .Y(n528) );
  OAI21XLTS U719 ( .A0(n529), .A1(n528), .B0(n1625), .Y(n527) );
  OAI31X1TS U720 ( .A0(n529), .A1(n1625), .A2(n528), .B0(n527), .Y(
        \mult_x_1/n960 ) );
  OAI22X1TS U721 ( .A0(n1602), .A1(n1401), .B0(n1601), .B1(n1460), .Y(n532) );
  OAI22X1TS U722 ( .A0(n927), .A1(n1492), .B0(n394), .B1(n1495), .Y(n531) );
  OAI21XLTS U723 ( .A0(n532), .A1(n531), .B0(n1671), .Y(n530) );
  OAI31X1TS U724 ( .A0(n532), .A1(n1671), .A2(n531), .B0(n530), .Y(
        \mult_x_1/n989 ) );
  OAI22X1TS U725 ( .A0(n723), .A1(n1561), .B0(n727), .B1(n1650), .Y(n535) );
  OAI22X1TS U726 ( .A0(n1643), .A1(n1580), .B0(n1642), .B1(n1560), .Y(n534) );
  OAI21XLTS U727 ( .A0(n535), .A1(n534), .B0(n1621), .Y(n533) );
  OAI31X1TS U728 ( .A0(n535), .A1(n1621), .A2(n534), .B0(n533), .Y(
        \mult_x_1/n1016 ) );
  OAI22X1TS U729 ( .A0(n723), .A1(n1440), .B0(n727), .B1(n1580), .Y(n538) );
  OAI22X1TS U730 ( .A0(n1643), .A1(n1560), .B0(n1642), .B1(n1454), .Y(n537) );
  OAI21XLTS U731 ( .A0(n538), .A1(n537), .B0(n1621), .Y(n536) );
  OAI31X1TS U732 ( .A0(n538), .A1(n1621), .A2(n537), .B0(n536), .Y(
        \mult_x_1/n1017 ) );
  INVX2TS U733 ( .A(A[18]), .Y(n542) );
  OAI22X1TS U734 ( .A0(n539), .A1(n542), .B0(A[18]), .B1(A[17]), .Y(n605) );
  INVX2TS U735 ( .A(n605), .Y(n985) );
  INVX2TS U736 ( .A(A[19]), .Y(n541) );
  OAI22X1TS U737 ( .A0(n1672), .A1(n541), .B0(A[19]), .B1(A[20]), .Y(n606) );
  INVX2TS U738 ( .A(n606), .Y(n543) );
  OAI22X1TS U739 ( .A0(n542), .A1(A[19]), .B0(n541), .B1(A[18]), .Y(n604) );
  INVX2TS U740 ( .A(n604), .Y(n544) );
  AND3X1TS U741 ( .A(n605), .B(n544), .C(n543), .Y(n986) );
  INVX2TS U742 ( .A(n986), .Y(n1003) );
  OAI22X1TS U743 ( .A0(n989), .A1(n1662), .B0(n1003), .B1(n1664), .Y(n545) );
  XOR2XLTS U744 ( .A(A[20]), .B(n545), .Y(\mult_x_1/n1048 ) );
  OAI22X1TS U745 ( .A0(n723), .A1(n1453), .B0(n727), .B1(n1560), .Y(n548) );
  OAI22X1TS U746 ( .A0(n1643), .A1(n1454), .B0(n1642), .B1(n1475), .Y(n547) );
  OAI21XLTS U747 ( .A0(n548), .A1(n547), .B0(n1621), .Y(n546) );
  OAI31X1TS U748 ( .A0(n548), .A1(n1621), .A2(n547), .B0(n546), .Y(
        \mult_x_1/n1018 ) );
  OAI22X1TS U749 ( .A0(n1565), .A1(n1444), .B0(n1564), .B1(n1470), .Y(n551) );
  OAI22X1TS U750 ( .A0(n319), .A1(n1479), .B0(n322), .B1(n1482), .Y(n550) );
  OAI21XLTS U751 ( .A0(n551), .A1(n550), .B0(A[29]), .Y(n549) );
  OAI31X1TS U752 ( .A0(n551), .A1(A[29]), .A2(n550), .B0(n549), .Y(n589) );
  NOR2XLTS U753 ( .A(n1468), .B(n1579), .Y(n553) );
  OAI22X1TS U754 ( .A0(n1414), .A1(n1592), .B0(n1413), .B1(n1559), .Y(n552) );
  AOI211XLTS U755 ( .A0(n1584), .A1(B[11]), .B0(n553), .C0(n552), .Y(n588) );
  INVX2TS U756 ( .A(n554), .Y(\mult_x_1/n426 ) );
  OAI22X1TS U757 ( .A0(n1602), .A1(n1427), .B0(n1601), .B1(n1461), .Y(n557) );
  OAI22X1TS U758 ( .A0(n927), .A1(n1460), .B0(n394), .B1(n1492), .Y(n556) );
  OAI21XLTS U759 ( .A0(n557), .A1(n556), .B0(n1671), .Y(n555) );
  OAI31X1TS U760 ( .A0(n557), .A1(n1671), .A2(n556), .B0(n555), .Y(
        \mult_x_1/n990 ) );
  OAI22X1TS U761 ( .A0(n1565), .A1(n1469), .B0(n1564), .B1(n1468), .Y(n560) );
  OAI22X1TS U762 ( .A0(n796), .A1(n1470), .B0(n322), .B1(n1479), .Y(n559) );
  OAI21XLTS U763 ( .A0(n560), .A1(n559), .B0(A[29]), .Y(n558) );
  OAI31X1TS U764 ( .A0(n560), .A1(A[29]), .A2(n559), .B0(n558), .Y(n586) );
  NOR2XLTS U765 ( .A(n1435), .B(n1579), .Y(n562) );
  OAI22X1TS U766 ( .A0(n1409), .A1(n1592), .B0(n1419), .B1(n1559), .Y(n561) );
  AOI211XLTS U767 ( .A0(n1584), .A1(B[10]), .B0(n562), .C0(n561), .Y(n585) );
  INVX2TS U768 ( .A(n563), .Y(\mult_x_1/n439 ) );
  OAI22X1TS U769 ( .A0(n723), .A1(n1397), .B0(n727), .B1(n1454), .Y(n566) );
  OAI22X1TS U770 ( .A0(n1643), .A1(n1475), .B0(n1642), .B1(n1487), .Y(n565) );
  OAI21XLTS U771 ( .A0(n566), .A1(n565), .B0(n1621), .Y(n564) );
  OAI31X1TS U772 ( .A0(n566), .A1(n1621), .A2(n565), .B0(n564), .Y(
        \mult_x_1/n1019 ) );
  INVX2TS U773 ( .A(\mult_x_1/n431 ), .Y(n596) );
  INVX2TS U774 ( .A(\mult_x_1/n419 ), .Y(n595) );
  INVX2TS U775 ( .A(n570), .Y(Product[42]) );
  INVX2TS U776 ( .A(n572), .Y(\mult_x_1/n493 ) );
  OAI22X1TS U777 ( .A0(n1565), .A1(n1436), .B0(n1564), .B1(n1435), .Y(n575) );
  OAI22X1TS U778 ( .A0(n319), .A1(n1468), .B0(n322), .B1(n1470), .Y(n574) );
  OAI21XLTS U779 ( .A0(n575), .A1(n574), .B0(n1625), .Y(n573) );
  OAI31X1TS U780 ( .A0(n575), .A1(n1625), .A2(n574), .B0(n573), .Y(
        \mult_x_1/n963 ) );
  OAI22X1TS U781 ( .A0(n1602), .A1(n1459), .B0(n1601), .B1(n1458), .Y(n578) );
  OAI22X1TS U782 ( .A0(n927), .A1(n1461), .B0(n394), .B1(n1460), .Y(n577) );
  OAI21XLTS U783 ( .A0(n578), .A1(n577), .B0(n1671), .Y(n576) );
  OAI31X1TS U784 ( .A0(n578), .A1(n1671), .A2(n577), .B0(n576), .Y(
        \mult_x_1/n991 ) );
  OAI22X1TS U785 ( .A0(n1602), .A1(n1393), .B0(n1601), .B1(n1449), .Y(n581) );
  OAI22X1TS U786 ( .A0(n927), .A1(n1458), .B0(n394), .B1(n1461), .Y(n580) );
  OAI21XLTS U787 ( .A0(n581), .A1(n580), .B0(n1671), .Y(n579) );
  OAI31X1TS U788 ( .A0(n581), .A1(n1671), .A2(n580), .B0(n579), .Y(
        \mult_x_1/n992 ) );
  OAI22X1TS U789 ( .A0(n723), .A1(n1474), .B0(n727), .B1(n1475), .Y(n584) );
  OAI22X1TS U790 ( .A0(n1643), .A1(n1487), .B0(n1642), .B1(n1488), .Y(n583) );
  OAI21XLTS U791 ( .A0(n584), .A1(n583), .B0(n1621), .Y(n582) );
  OAI31X1TS U792 ( .A0(n584), .A1(n1621), .A2(n583), .B0(n582), .Y(
        \mult_x_1/n1020 ) );
  INVX2TS U793 ( .A(n587), .Y(\mult_x_1/n440 ) );
  INVX2TS U794 ( .A(n590), .Y(\mult_x_1/n427 ) );
  OAI22X1TS U795 ( .A0(n723), .A1(n1486), .B0(n727), .B1(n1487), .Y(n593) );
  OAI22X1TS U796 ( .A0(n1643), .A1(n1488), .B0(n1640), .B1(n1494), .Y(n592) );
  OAI21XLTS U797 ( .A0(n593), .A1(n592), .B0(n1621), .Y(n591) );
  OAI31X1TS U798 ( .A0(n593), .A1(n1621), .A2(n592), .B0(n591), .Y(
        \mult_x_1/n1021 ) );
  INVX2TS U799 ( .A(\mult_x_1/n418 ), .Y(n651) );
  INVX2TS U800 ( .A(\mult_x_1/n408 ), .Y(n650) );
  INVX2TS U801 ( .A(n597), .Y(Product[43]) );
  OAI22X1TS U802 ( .A0(n1565), .A1(n1409), .B0(n1564), .B1(n1419), .Y(n600) );
  OAI22X1TS U803 ( .A0(n319), .A1(n1413), .B0(n322), .B1(n1435), .Y(n599) );
  OAI21XLTS U804 ( .A0(n600), .A1(n599), .B0(n1625), .Y(n598) );
  OAI31X1TS U805 ( .A0(n600), .A1(n1625), .A2(n599), .B0(n598), .Y(
        \mult_x_1/n965 ) );
  OAI22X1TS U806 ( .A0(n1565), .A1(n1414), .B0(n1564), .B1(n1413), .Y(n603) );
  OAI22X1TS U807 ( .A0(n319), .A1(n1435), .B0(n322), .B1(n1468), .Y(n602) );
  OAI21XLTS U808 ( .A0(n603), .A1(n602), .B0(n1625), .Y(n601) );
  OAI31X1TS U809 ( .A0(n603), .A1(n1625), .A2(n602), .B0(n601), .Y(
        \mult_x_1/n964 ) );
  OAI22X1TS U810 ( .A0(n989), .A1(n1581), .B0(n1003), .B1(n1580), .Y(n609) );
  CLKAND2X2TS U811 ( .A(n605), .B(n604), .Y(n991) );
  CLKAND2X2TS U812 ( .A(n606), .B(n985), .Y(n987) );
  INVX2TS U813 ( .A(n987), .Y(n1005) );
  OAI22X1TS U814 ( .A0(n1004), .A1(n1650), .B0(n1005), .B1(n1664), .Y(n608) );
  OAI21XLTS U815 ( .A0(n609), .A1(n608), .B0(n1672), .Y(n607) );
  OAI31X1TS U816 ( .A0(n609), .A1(n1672), .A2(n608), .B0(n607), .Y(
        \mult_x_1/n1050 ) );
  OAI22X1TS U817 ( .A0(n1602), .A1(n1448), .B0(n1601), .B1(n1482), .Y(n612) );
  OAI22X1TS U818 ( .A0(n927), .A1(n1481), .B0(n394), .B1(n1449), .Y(n611) );
  OAI21XLTS U819 ( .A0(n612), .A1(n611), .B0(n1671), .Y(n610) );
  OAI31X1TS U820 ( .A0(n612), .A1(n1671), .A2(n611), .B0(n610), .Y(
        \mult_x_1/n994 ) );
  OAI22X1TS U821 ( .A0(n1602), .A1(n1423), .B0(n1601), .B1(n1481), .Y(n615) );
  OAI22X1TS U822 ( .A0(n927), .A1(n1449), .B0(n394), .B1(n1458), .Y(n614) );
  OAI21XLTS U823 ( .A0(n615), .A1(n614), .B0(n1671), .Y(n613) );
  OAI31X1TS U824 ( .A0(n615), .A1(n1671), .A2(n614), .B0(n613), .Y(
        \mult_x_1/n993 ) );
  OAI22X1TS U825 ( .A0(n1565), .A1(n1405), .B0(n1564), .B1(n1501), .Y(n618) );
  OAI22X1TS U826 ( .A0(n319), .A1(n1419), .B0(n322), .B1(n1413), .Y(n617) );
  OAI21XLTS U827 ( .A0(n618), .A1(n617), .B0(n1625), .Y(n616) );
  OAI31X1TS U828 ( .A0(n618), .A1(n1625), .A2(n617), .B0(n616), .Y(
        \mult_x_1/n966 ) );
  OAI22X1TS U829 ( .A0(n723), .A1(n1493), .B0(n727), .B1(n1494), .Y(n621) );
  OAI22X1TS U830 ( .A0(n1643), .A1(n1495), .B0(n1640), .B1(n1492), .Y(n620) );
  OAI21XLTS U831 ( .A0(n621), .A1(n620), .B0(n1621), .Y(n619) );
  OAI31X1TS U832 ( .A0(n621), .A1(n1621), .A2(n620), .B0(n619), .Y(
        \mult_x_1/n1023 ) );
  OAI22X1TS U833 ( .A0(n723), .A1(n1431), .B0(n727), .B1(n1488), .Y(n624) );
  OAI22X1TS U834 ( .A0(n1643), .A1(n1494), .B0(n1640), .B1(n1495), .Y(n623) );
  OAI21XLTS U835 ( .A0(n624), .A1(n623), .B0(n1621), .Y(n622) );
  OAI31X1TS U836 ( .A0(n624), .A1(n1621), .A2(n623), .B0(n622), .Y(
        \mult_x_1/n1022 ) );
  OAI22X1TS U837 ( .A0(n1602), .A1(n1480), .B0(n1601), .B1(n1479), .Y(n627) );
  OAI22X1TS U838 ( .A0(n927), .A1(n1482), .B0(n394), .B1(n1481), .Y(n626) );
  OAI21XLTS U839 ( .A0(n627), .A1(n626), .B0(n1671), .Y(n625) );
  OAI31X1TS U840 ( .A0(n627), .A1(n1671), .A2(n626), .B0(n625), .Y(
        \mult_x_1/n995 ) );
  OAI22X1TS U841 ( .A0(n1602), .A1(n1469), .B0(n1601), .B1(n1468), .Y(n630) );
  OAI22X1TS U842 ( .A0(n927), .A1(n1470), .B0(n394), .B1(n1479), .Y(n629) );
  OAI21XLTS U843 ( .A0(n630), .A1(n629), .B0(n1671), .Y(n628) );
  OAI31X1TS U844 ( .A0(n630), .A1(n1671), .A2(n629), .B0(n628), .Y(
        \mult_x_1/n997 ) );
  OAI22X1TS U845 ( .A0(n1602), .A1(n1444), .B0(n1601), .B1(n1470), .Y(n633) );
  OAI22X1TS U846 ( .A0(n927), .A1(n1479), .B0(n394), .B1(n1482), .Y(n632) );
  OAI21XLTS U847 ( .A0(n633), .A1(n632), .B0(n1671), .Y(n631) );
  OAI31X1TS U848 ( .A0(n633), .A1(n1671), .A2(n632), .B0(n631), .Y(
        \mult_x_1/n996 ) );
  OAI22X1TS U849 ( .A0(n723), .A1(n1401), .B0(n727), .B1(n1495), .Y(n636) );
  OAI22X1TS U850 ( .A0(n1643), .A1(n1492), .B0(n1640), .B1(n1460), .Y(n635) );
  OAI21XLTS U851 ( .A0(n636), .A1(n635), .B0(n1621), .Y(n634) );
  OAI31X1TS U852 ( .A0(n636), .A1(n1621), .A2(n635), .B0(n634), .Y(
        \mult_x_1/n1024 ) );
  OAI22X1TS U853 ( .A0(n989), .A1(n1561), .B0(n1003), .B1(n1560), .Y(n639) );
  OAI22X1TS U854 ( .A0(n1004), .A1(n1580), .B0(n1005), .B1(n1650), .Y(n638) );
  OAI21XLTS U855 ( .A0(n639), .A1(n638), .B0(n1672), .Y(n637) );
  OAI31X1TS U856 ( .A0(n639), .A1(n1672), .A2(n638), .B0(n637), .Y(
        \mult_x_1/n1051 ) );
  OAI22X1TS U857 ( .A0(n989), .A1(n1440), .B0(n1003), .B1(n1454), .Y(n642) );
  INVX2TS U858 ( .A(n991), .Y(n1004) );
  OAI22X1TS U859 ( .A0(n1004), .A1(n1560), .B0(n1005), .B1(n1580), .Y(n641) );
  OAI21XLTS U860 ( .A0(n642), .A1(n641), .B0(n1672), .Y(n640) );
  OAI31X1TS U861 ( .A0(n642), .A1(n1672), .A2(n641), .B0(n640), .Y(
        \mult_x_1/n1052 ) );
  OAI22X1TS U862 ( .A0(n1565), .A1(n1500), .B0(n1564), .B1(n1533), .Y(n645) );
  OAI22X1TS U863 ( .A0(n319), .A1(n1506), .B0(n322), .B1(n1501), .Y(n644) );
  OAI21XLTS U864 ( .A0(n645), .A1(n644), .B0(A[29]), .Y(n643) );
  OAI31X1TS U865 ( .A0(n645), .A1(A[29]), .A2(n644), .B0(n643), .Y(n689) );
  NOR2XLTS U866 ( .A(n1552), .B(n1579), .Y(n647) );
  OAI22X1TS U867 ( .A0(n1554), .A1(n1559), .B0(n1553), .B1(n1592), .Y(n646) );
  AOI211XLTS U868 ( .A0(n1584), .A1(B[4]), .B0(n647), .C0(n646), .Y(n688) );
  INVX2TS U869 ( .A(n648), .Y(\mult_x_1/n520 ) );
  INVX2TS U870 ( .A(\mult_x_1/n407 ), .Y(n677) );
  INVX2TS U871 ( .A(\mult_x_1/n398 ), .Y(n676) );
  INVX2TS U872 ( .A(n652), .Y(Product[44]) );
  INVX2TS U873 ( .A(n540), .Y(n989) );
  OAI22X1TS U874 ( .A0(n989), .A1(n1453), .B0(n1003), .B1(n1475), .Y(n655) );
  OAI22X1TS U875 ( .A0(n1004), .A1(n1454), .B0(n1005), .B1(n1560), .Y(n654) );
  OAI21XLTS U876 ( .A0(n655), .A1(n654), .B0(n1672), .Y(n653) );
  OAI31X1TS U877 ( .A0(n655), .A1(n1672), .A2(n654), .B0(n653), .Y(
        \mult_x_1/n1053 ) );
  AOI222XLTS U878 ( .A0(n540), .A1(n1606), .B0(n991), .B1(B[31]), .C0(n986), 
        .C1(B[30]), .Y(n656) );
  XOR2XLTS U879 ( .A(n1672), .B(n656), .Y(\mult_x_1/n1049 ) );
  OAI22X1TS U880 ( .A0(n1565), .A1(n1505), .B0(n1564), .B1(n1552), .Y(n659) );
  OAI22X1TS U881 ( .A0(n319), .A1(n1533), .B0(n322), .B1(n1506), .Y(n658) );
  OAI21XLTS U882 ( .A0(n659), .A1(n658), .B0(A[29]), .Y(n657) );
  OAI31X1TS U883 ( .A0(n659), .A1(A[29]), .A2(n658), .B0(n657), .Y(n692) );
  NOR2XLTS U884 ( .A(n813), .B(n1579), .Y(n661) );
  OAI22X1TS U885 ( .A0(n29), .A1(n1559), .B0(n1537), .B1(n1592), .Y(n660) );
  AOI211XLTS U886 ( .A0(n1584), .A1(B[3]), .B0(n661), .C0(n660), .Y(n691) );
  INVX2TS U887 ( .A(n662), .Y(\mult_x_1/n534 ) );
  OAI22X1TS U888 ( .A0(n1565), .A1(n1418), .B0(n1564), .B1(n1506), .Y(n665) );
  OAI22X1TS U889 ( .A0(n319), .A1(n1501), .B0(n322), .B1(n1419), .Y(n664) );
  OAI21XLTS U890 ( .A0(n665), .A1(n664), .B0(A[29]), .Y(n663) );
  OAI31X1TS U891 ( .A0(n665), .A1(A[29]), .A2(n664), .B0(n663), .Y(n686) );
  NOR2XLTS U892 ( .A(n1533), .B(n1579), .Y(n667) );
  OAI22X1TS U893 ( .A0(n1532), .A1(n1592), .B0(n813), .B1(n1559), .Y(n666) );
  AOI211XLTS U894 ( .A0(n1584), .A1(B[5]), .B0(n667), .C0(n666), .Y(n685) );
  INVX2TS U895 ( .A(n668), .Y(\mult_x_1/n506 ) );
  OAI22X1TS U896 ( .A0(n723), .A1(n1427), .B0(n727), .B1(n1492), .Y(n671) );
  OAI22X1TS U897 ( .A0(n1643), .A1(n1460), .B0(n1640), .B1(n1461), .Y(n670) );
  OAI21XLTS U898 ( .A0(n671), .A1(n670), .B0(n1621), .Y(n669) );
  OAI31X1TS U899 ( .A0(n671), .A1(n1621), .A2(n670), .B0(n669), .Y(
        \mult_x_1/n1025 ) );
  OAI22X1TS U900 ( .A0(n989), .A1(n1397), .B0(n1003), .B1(n1487), .Y(n674) );
  OAI22X1TS U901 ( .A0(n1004), .A1(n1475), .B0(n1005), .B1(n1454), .Y(n673) );
  OAI21XLTS U902 ( .A0(n674), .A1(n673), .B0(n1672), .Y(n672) );
  OAI31X1TS U903 ( .A0(n674), .A1(n1672), .A2(n673), .B0(n672), .Y(
        \mult_x_1/n1054 ) );
  INVX2TS U904 ( .A(\mult_x_1/n397 ), .Y(n715) );
  INVX2TS U905 ( .A(\mult_x_1/n387 ), .Y(n714) );
  INVX2TS U906 ( .A(n678), .Y(Product[45]) );
  OAI22X1TS U907 ( .A0(n1602), .A1(n1436), .B0(n1601), .B1(n1435), .Y(n681) );
  OAI22X1TS U908 ( .A0(n927), .A1(n1468), .B0(n394), .B1(n1470), .Y(n680) );
  OAI21XLTS U909 ( .A0(n681), .A1(n680), .B0(n1671), .Y(n679) );
  OAI31X1TS U910 ( .A0(n681), .A1(n1671), .A2(n680), .B0(n679), .Y(
        \mult_x_1/n998 ) );
  OAI22X1TS U911 ( .A0(n723), .A1(n1459), .B0(n727), .B1(n1460), .Y(n684) );
  OAI22X1TS U912 ( .A0(n1643), .A1(n1461), .B0(n1640), .B1(n1458), .Y(n683) );
  OAI21XLTS U913 ( .A0(n684), .A1(n683), .B0(n1621), .Y(n682) );
  OAI31X1TS U914 ( .A0(n684), .A1(n1621), .A2(n683), .B0(n682), .Y(
        \mult_x_1/n1026 ) );
  INVX2TS U915 ( .A(n687), .Y(\mult_x_1/n507 ) );
  INVX2TS U916 ( .A(n690), .Y(\mult_x_1/n521 ) );
  INVX2TS U917 ( .A(n694), .Y(\mult_x_1/n535 ) );
  OAI22X1TS U918 ( .A0(n723), .A1(n1393), .B0(n727), .B1(n1461), .Y(n697) );
  OAI22X1TS U919 ( .A0(n1643), .A1(n1458), .B0(n1640), .B1(n1449), .Y(n696) );
  OAI21XLTS U920 ( .A0(n697), .A1(n696), .B0(n1621), .Y(n695) );
  OAI31X1TS U921 ( .A0(n697), .A1(n1621), .A2(n696), .B0(n695), .Y(
        \mult_x_1/n1027 ) );
  OAI22X1TS U922 ( .A0(n989), .A1(n1474), .B0(n1003), .B1(n1488), .Y(n700) );
  OAI22X1TS U923 ( .A0(n1004), .A1(n1487), .B0(n1005), .B1(n1475), .Y(n699) );
  OAI21XLTS U924 ( .A0(n700), .A1(n699), .B0(n1672), .Y(n698) );
  OAI31X1TS U925 ( .A0(n700), .A1(n1672), .A2(n699), .B0(n698), .Y(
        \mult_x_1/n1055 ) );
  OAI22X1TS U926 ( .A0(n989), .A1(n1486), .B0(n1003), .B1(n1494), .Y(n703) );
  OAI22X1TS U927 ( .A0(n1004), .A1(n1488), .B0(n1005), .B1(n1487), .Y(n702) );
  OAI21XLTS U928 ( .A0(n703), .A1(n702), .B0(n1672), .Y(n701) );
  OAI31X1TS U929 ( .A0(n703), .A1(n1672), .A2(n702), .B0(n701), .Y(
        \mult_x_1/n1056 ) );
  OAI22X1TS U930 ( .A0(n1602), .A1(n1409), .B0(n1601), .B1(n1419), .Y(n706) );
  INVX2TS U931 ( .A(n899), .Y(n902) );
  OAI22X1TS U932 ( .A0(n927), .A1(n1413), .B0(n902), .B1(n1435), .Y(n705) );
  OAI21XLTS U933 ( .A0(n706), .A1(n705), .B0(n1671), .Y(n704) );
  OAI31X1TS U934 ( .A0(n706), .A1(n1671), .A2(n705), .B0(n704), .Y(
        \mult_x_1/n1000 ) );
  OAI22X1TS U935 ( .A0(n1602), .A1(n1405), .B0(n1601), .B1(n1501), .Y(n709) );
  OAI22X1TS U936 ( .A0(n927), .A1(n1419), .B0(n902), .B1(n1413), .Y(n708) );
  OAI21XLTS U937 ( .A0(n709), .A1(n708), .B0(n1671), .Y(n707) );
  OAI31X1TS U938 ( .A0(n709), .A1(n1671), .A2(n708), .B0(n707), .Y(
        \mult_x_1/n1001 ) );
  OAI22X1TS U939 ( .A0(n1602), .A1(n1414), .B0(n1601), .B1(n1413), .Y(n712) );
  OAI22X1TS U940 ( .A0(n927), .A1(n1435), .B0(n394), .B1(n1468), .Y(n711) );
  OAI21XLTS U941 ( .A0(n712), .A1(n711), .B0(n1671), .Y(n710) );
  OAI31X1TS U942 ( .A0(n712), .A1(n1671), .A2(n711), .B0(n710), .Y(
        \mult_x_1/n999 ) );
  INVX2TS U943 ( .A(\mult_x_1/n386 ), .Y(n739) );
  INVX2TS U944 ( .A(\mult_x_1/n379 ), .Y(n738) );
  INVX2TS U945 ( .A(n716), .Y(Product[46]) );
  OAI2BB2XLTS U946 ( .B0(n1673), .B1(A[15]), .A0N(A[15]), .A1N(n1673), .Y(n719) );
  INVX2TS U947 ( .A(n719), .Y(n1263) );
  OAI2BB2XLTS U948 ( .B0(A[16]), .B1(A[17]), .A0N(A[17]), .A1N(A[16]), .Y(n718) );
  NOR2XLTS U949 ( .A(n1263), .B(n718), .Y(n1607) );
  INVX2TS U950 ( .A(n1607), .Y(n1646) );
  XOR2XLTS U951 ( .A(A[15]), .B(A[16]), .Y(n717) );
  NOR3XLTS U952 ( .A(n718), .B(n719), .C(n717), .Y(n1604) );
  INVX2TS U953 ( .A(n1604), .Y(n1645) );
  OAI22X1TS U954 ( .A0(n1646), .A1(n1581), .B0(n1645), .B1(n1580), .Y(n722) );
  NAND2X1TS U955 ( .A(n717), .B(n1263), .Y(n1346) );
  INVX2TS U956 ( .A(n1346), .Y(n1605) );
  INVX2TS U957 ( .A(n1605), .Y(n1361) );
  OAI22X1TS U958 ( .A0(n1361), .A1(n1650), .B0(n1264), .B1(n1664), .Y(n721) );
  OAI21XLTS U959 ( .A0(n722), .A1(n721), .B0(n539), .Y(n720) );
  OAI31X1TS U960 ( .A0(n722), .A1(n539), .A2(n721), .B0(n720), .Y(
        \mult_x_1/n1085 ) );
  OAI22X1TS U961 ( .A0(n723), .A1(n1423), .B0(n727), .B1(n1458), .Y(n726) );
  OAI22X1TS U962 ( .A0(n1643), .A1(n1449), .B0(n1640), .B1(n1481), .Y(n725) );
  OAI21XLTS U963 ( .A0(n726), .A1(n725), .B0(n1621), .Y(n724) );
  OAI31X1TS U964 ( .A0(n726), .A1(n1621), .A2(n725), .B0(n724), .Y(
        \mult_x_1/n1028 ) );
  OAI22X1TS U965 ( .A0(n723), .A1(n1448), .B0(n727), .B1(n1449), .Y(n730) );
  OAI22X1TS U966 ( .A0(n1643), .A1(n1481), .B0(n1640), .B1(n1482), .Y(n729) );
  OAI21XLTS U967 ( .A0(n730), .A1(n729), .B0(n1621), .Y(n728) );
  OAI31X1TS U968 ( .A0(n730), .A1(n1621), .A2(n729), .B0(n728), .Y(
        \mult_x_1/n1029 ) );
  OAI22X1TS U969 ( .A0(n1602), .A1(n1418), .B0(n1601), .B1(n1506), .Y(n733) );
  OAI22X1TS U970 ( .A0(n927), .A1(n1501), .B0(n902), .B1(n1419), .Y(n732) );
  OAI21XLTS U971 ( .A0(n733), .A1(n732), .B0(n1671), .Y(n731) );
  OAI31X1TS U972 ( .A0(n733), .A1(n1671), .A2(n732), .B0(n731), .Y(
        \mult_x_1/n1002 ) );
  OAI22X1TS U973 ( .A0(n1602), .A1(n1500), .B0(n1601), .B1(n1533), .Y(n736) );
  OAI22X1TS U974 ( .A0(n927), .A1(n1506), .B0(n902), .B1(n1501), .Y(n735) );
  OAI21XLTS U975 ( .A0(n736), .A1(n735), .B0(n1671), .Y(n734) );
  OAI31X1TS U976 ( .A0(n736), .A1(n1671), .A2(n735), .B0(n734), .Y(
        \mult_x_1/n1003 ) );
  INVX2TS U977 ( .A(\mult_x_1/n378 ), .Y(n819) );
  INVX2TS U978 ( .A(\mult_x_1/n370 ), .Y(n818) );
  INVX2TS U979 ( .A(n740), .Y(Product[47]) );
  OAI22X1TS U980 ( .A0(n989), .A1(n1493), .B0(n1003), .B1(n1492), .Y(n743) );
  OAI22X1TS U981 ( .A0(n1004), .A1(n1495), .B0(n1005), .B1(n1494), .Y(n742) );
  OAI21XLTS U982 ( .A0(n743), .A1(n742), .B0(n1672), .Y(n741) );
  OAI31X1TS U983 ( .A0(n743), .A1(n1672), .A2(n742), .B0(n741), .Y(
        \mult_x_1/n1058 ) );
  OAI22X1TS U984 ( .A0(n989), .A1(n1431), .B0(n1003), .B1(n1495), .Y(n746) );
  OAI22X1TS U985 ( .A0(n1004), .A1(n1494), .B0(n1005), .B1(n1488), .Y(n745) );
  OAI21XLTS U986 ( .A0(n746), .A1(n745), .B0(n1672), .Y(n744) );
  OAI31X1TS U987 ( .A0(n746), .A1(n1672), .A2(n745), .B0(n744), .Y(
        \mult_x_1/n1057 ) );
  OAI22X1TS U988 ( .A0(n723), .A1(n1480), .B0(n727), .B1(n1481), .Y(n749) );
  OAI22X1TS U989 ( .A0(n1643), .A1(n1482), .B0(n1640), .B1(n1479), .Y(n748) );
  OAI21XLTS U990 ( .A0(n749), .A1(n748), .B0(n1621), .Y(n747) );
  OAI31X1TS U991 ( .A0(n749), .A1(n1621), .A2(n748), .B0(n747), .Y(
        \mult_x_1/n1030 ) );
  OAI22X1TS U992 ( .A0(n1602), .A1(n1505), .B0(n1601), .B1(n1552), .Y(n752) );
  OAI22X1TS U993 ( .A0(n927), .A1(n1533), .B0(n394), .B1(n1506), .Y(n751) );
  OAI21XLTS U994 ( .A0(n752), .A1(n751), .B0(n1671), .Y(n750) );
  OAI31X1TS U995 ( .A0(n752), .A1(n1671), .A2(n751), .B0(n750), .Y(
        \mult_x_1/n1004 ) );
  OAI22X1TS U996 ( .A0(n723), .A1(n1444), .B0(n727), .B1(n1482), .Y(n755) );
  OAI22X1TS U997 ( .A0(n1643), .A1(n1479), .B0(n1640), .B1(n1470), .Y(n754) );
  OAI21XLTS U998 ( .A0(n755), .A1(n754), .B0(n1621), .Y(n753) );
  OAI31X1TS U999 ( .A0(n755), .A1(n1621), .A2(n754), .B0(n753), .Y(
        \mult_x_1/n1031 ) );
  OAI22X1TS U1000 ( .A0(n723), .A1(n1469), .B0(n727), .B1(n1479), .Y(n758) );
  OAI22X1TS U1001 ( .A0(n1643), .A1(n1470), .B0(n1640), .B1(n1468), .Y(n757)
         );
  OAI21XLTS U1002 ( .A0(n758), .A1(n757), .B0(n1621), .Y(n756) );
  OAI31X1TS U1003 ( .A0(n758), .A1(n1621), .A2(n757), .B0(n756), .Y(
        \mult_x_1/n1032 ) );
  OAI22X1TS U1004 ( .A0(n989), .A1(n1401), .B0(n1003), .B1(n1460), .Y(n761) );
  OAI22X1TS U1005 ( .A0(n1004), .A1(n1492), .B0(n1005), .B1(n1495), .Y(n760)
         );
  OAI21XLTS U1006 ( .A0(n761), .A1(n760), .B0(n1672), .Y(n759) );
  OAI31X1TS U1007 ( .A0(n761), .A1(n1672), .A2(n760), .B0(n759), .Y(
        \mult_x_1/n1059 ) );
  OAI22X1TS U1008 ( .A0(n1646), .A1(n1561), .B0(n1645), .B1(n1560), .Y(n764)
         );
  OAI22X1TS U1009 ( .A0(n1361), .A1(n1580), .B0(n1264), .B1(n1650), .Y(n763)
         );
  OAI21XLTS U1010 ( .A0(n764), .A1(n763), .B0(n539), .Y(n762) );
  OAI31X1TS U1011 ( .A0(n764), .A1(n539), .A2(n763), .B0(n762), .Y(
        \mult_x_1/n1086 ) );
  OAI22X1TS U1012 ( .A0(n1646), .A1(n1440), .B0(n1645), .B1(n1454), .Y(n767)
         );
  OAI22X1TS U1013 ( .A0(n1361), .A1(n1560), .B0(n1264), .B1(n1580), .Y(n766)
         );
  OAI21XLTS U1014 ( .A0(n767), .A1(n766), .B0(n539), .Y(n765) );
  OAI31X1TS U1015 ( .A0(n767), .A1(n539), .A2(n766), .B0(n765), .Y(
        \mult_x_1/n1087 ) );
  INVX2TS U1016 ( .A(A[12]), .Y(n769) );
  OAI22X1TS U1017 ( .A0(n1638), .A1(n769), .B0(A[12]), .B1(A[11]), .Y(n857) );
  INVX2TS U1018 ( .A(n857), .Y(n1181) );
  INVX2TS U1019 ( .A(A[13]), .Y(n768) );
  OAI22X1TS U1020 ( .A0(n1673), .A1(n768), .B0(A[13]), .B1(A[14]), .Y(n858) );
  INVX2TS U1021 ( .A(n858), .Y(n770) );
  CLKAND2X2TS U1022 ( .A(n1181), .B(n770), .Y(n1182) );
  INVX2TS U1023 ( .A(n1182), .Y(n1186) );
  OAI22X1TS U1024 ( .A0(n769), .A1(A[13]), .B0(n768), .B1(A[12]), .Y(n856) );
  INVX2TS U1025 ( .A(n856), .Y(n771) );
  INVX2TS U1026 ( .A(n1), .Y(n1175) );
  OAI22X1TS U1027 ( .A0(n1186), .A1(n1662), .B0(n1175), .B1(n1664), .Y(n772)
         );
  XOR2XLTS U1028 ( .A(A[14]), .B(n772), .Y(\mult_x_1/n1118 ) );
  OAI22X1TS U1029 ( .A0(n1646), .A1(n1453), .B0(n1645), .B1(n1475), .Y(n775)
         );
  OAI22X1TS U1030 ( .A0(n1361), .A1(n1454), .B0(n1264), .B1(n1560), .Y(n774)
         );
  OAI21XLTS U1031 ( .A0(n775), .A1(n774), .B0(n539), .Y(n773) );
  OAI31X1TS U1032 ( .A0(n775), .A1(n539), .A2(n774), .B0(n773), .Y(
        \mult_x_1/n1088 ) );
  OAI22X1TS U1033 ( .A0(n1565), .A1(n1532), .B0(n1564), .B1(n813), .Y(n778) );
  OAI22X1TS U1034 ( .A0(n319), .A1(n1552), .B0(n322), .B1(n1533), .Y(n777) );
  OAI21XLTS U1035 ( .A0(n778), .A1(n777), .B0(A[29]), .Y(n776) );
  OAI31X1TS U1036 ( .A0(n778), .A1(A[29]), .A2(n777), .B0(n776), .Y(n836) );
  NOR2XLTS U1037 ( .A(n1554), .B(n1579), .Y(n780) );
  OAI22X1TS U1038 ( .A0(n1527), .A1(n1592), .B0(n23), .B1(n1559), .Y(n779) );
  AOI211XLTS U1039 ( .A0(n1584), .A1(B[2]), .B0(n780), .C0(n779), .Y(n835) );
  OAI22X1TS U1040 ( .A0(n1554), .A1(n1564), .B0(n1565), .B1(n1553), .Y(n783)
         );
  OAI22X1TS U1041 ( .A0(n319), .A1(n813), .B0(n322), .B1(n1552), .Y(n782) );
  OAI21XLTS U1042 ( .A0(n783), .A1(n782), .B0(A[29]), .Y(n781) );
  OAI31X1TS U1043 ( .A0(n783), .A1(A[29]), .A2(n782), .B0(n781), .Y(n847) );
  NOR2XLTS U1044 ( .A(n29), .B(n1579), .Y(n785) );
  OAI22X1TS U1045 ( .A0(n9), .A1(n1559), .B0(n1517), .B1(n1592), .Y(n784) );
  AOI211XLTS U1046 ( .A0(n1584), .A1(B[1]), .B0(n785), .C0(n784), .Y(n846) );
  OAI22X1TS U1047 ( .A0(n29), .A1(n1564), .B0(n1565), .B1(n1537), .Y(n788) );
  OAI22X1TS U1048 ( .A0(n1554), .A1(n796), .B0(n322), .B1(n813), .Y(n787) );
  OAI21XLTS U1049 ( .A0(n788), .A1(n787), .B0(A[29]), .Y(n786) );
  OAI31X1TS U1050 ( .A0(n788), .A1(A[29]), .A2(n787), .B0(n786), .Y(n843) );
  OAI222X1TS U1051 ( .A0(n23), .A1(n1579), .B0(n9), .B1(n1591), .C0(n1516), 
        .C1(n1592), .Y(n789) );
  INVX2TS U1052 ( .A(n789), .Y(n842) );
  NOR2XLTS U1053 ( .A(n9), .B(n790), .Y(\mult_x_1/n633 ) );
  OAI222X1TS U1054 ( .A0(n1565), .A1(n1516), .B0(n322), .B1(n23), .C0(n796), 
        .C1(n9), .Y(n852) );
  AOI21X1TS U1055 ( .A0(A[29]), .A1(\mult_x_1/n633 ), .B0(n852), .Y(n1623) );
  INVX2TS U1056 ( .A(n1623), .Y(n794) );
  OAI22X1TS U1057 ( .A0(n9), .A1(n1564), .B0(n1517), .B1(n1565), .Y(n792) );
  OAI22X1TS U1058 ( .A0(n29), .A1(n322), .B0(n23), .B1(n796), .Y(n791) );
  NOR2XLTS U1059 ( .A(n792), .B(n791), .Y(n1626) );
  NAND2X1TS U1060 ( .A(A[29]), .B(n1626), .Y(n793) );
  OR2X1TS U1061 ( .A(n794), .B(n793), .Y(n1622) );
  NAND2X1TS U1062 ( .A(B[0]), .B(n795), .Y(n840) );
  OAI22X1TS U1063 ( .A0(n1527), .A1(n1565), .B0(n23), .B1(n1564), .Y(n799) );
  OAI22X1TS U1064 ( .A0(n1554), .A1(n322), .B0(n29), .B1(n796), .Y(n798) );
  OAI21XLTS U1065 ( .A0(n799), .A1(n798), .B0(A[29]), .Y(n797) );
  OAI31X1TS U1066 ( .A0(n799), .A1(A[29]), .A2(n798), .B0(n797), .Y(n838) );
  AO21XLTS U1067 ( .A0(n1622), .A1(n840), .B0(n838), .Y(n841) );
  INVX2TS U1068 ( .A(n800), .Y(\mult_x_1/n548 ) );
  OAI22X1TS U1069 ( .A0(n989), .A1(n1427), .B0(n1003), .B1(n1461), .Y(n803) );
  OAI22X1TS U1070 ( .A0(n1004), .A1(n1460), .B0(n1005), .B1(n1492), .Y(n802)
         );
  OAI21XLTS U1071 ( .A0(n803), .A1(n802), .B0(n1672), .Y(n801) );
  OAI31X1TS U1072 ( .A0(n803), .A1(n1672), .A2(n802), .B0(n801), .Y(
        \mult_x_1/n1060 ) );
  OAI22X1TS U1073 ( .A0(n989), .A1(n1459), .B0(n1003), .B1(n1458), .Y(n806) );
  OAI22X1TS U1074 ( .A0(n1004), .A1(n1461), .B0(n1005), .B1(n1460), .Y(n805)
         );
  OAI21XLTS U1075 ( .A0(n806), .A1(n805), .B0(n1672), .Y(n804) );
  OAI31X1TS U1076 ( .A0(n806), .A1(n1672), .A2(n805), .B0(n804), .Y(
        \mult_x_1/n1061 ) );
  OAI22X1TS U1077 ( .A0(n1646), .A1(n1397), .B0(n1645), .B1(n1487), .Y(n809)
         );
  OAI22X1TS U1078 ( .A0(n1361), .A1(n1475), .B0(n1264), .B1(n1454), .Y(n808)
         );
  OAI21XLTS U1079 ( .A0(n809), .A1(n808), .B0(n539), .Y(n807) );
  OAI31X1TS U1080 ( .A0(n809), .A1(n539), .A2(n808), .B0(n807), .Y(
        \mult_x_1/n1089 ) );
  OAI22X1TS U1081 ( .A0(n723), .A1(n1436), .B0(n727), .B1(n1470), .Y(n812) );
  OAI22X1TS U1082 ( .A0(n1643), .A1(n1468), .B0(n1640), .B1(n1435), .Y(n811)
         );
  OAI21XLTS U1083 ( .A0(n812), .A1(n811), .B0(n1621), .Y(n810) );
  OAI31X1TS U1084 ( .A0(n812), .A1(n1621), .A2(n811), .B0(n810), .Y(
        \mult_x_1/n1033 ) );
  OAI22X1TS U1085 ( .A0(n1602), .A1(n1532), .B0(n1601), .B1(n813), .Y(n816) );
  OAI22X1TS U1086 ( .A0(n927), .A1(n1552), .B0(n902), .B1(n1533), .Y(n815) );
  OAI21XLTS U1087 ( .A0(n816), .A1(n815), .B0(n1671), .Y(n814) );
  OAI31X1TS U1088 ( .A0(n816), .A1(n1671), .A2(n815), .B0(n814), .Y(
        \mult_x_1/n1005 ) );
  INVX2TS U1089 ( .A(\mult_x_1/n369 ), .Y(n832) );
  INVX2TS U1090 ( .A(\mult_x_1/n360 ), .Y(n831) );
  INVX2TS U1091 ( .A(n820), .Y(Product[48]) );
  OAI22X1TS U1092 ( .A0(n989), .A1(n1393), .B0(n1003), .B1(n1449), .Y(n823) );
  OAI22X1TS U1093 ( .A0(n1004), .A1(n1458), .B0(n1005), .B1(n1461), .Y(n822)
         );
  OAI21XLTS U1094 ( .A0(n823), .A1(n822), .B0(n1672), .Y(n821) );
  OAI31X1TS U1095 ( .A0(n823), .A1(n1672), .A2(n822), .B0(n821), .Y(
        \mult_x_1/n1062 ) );
  OAI22X1TS U1096 ( .A0(n1646), .A1(n1474), .B0(n1645), .B1(n1488), .Y(n826)
         );
  OAI22X1TS U1097 ( .A0(n1361), .A1(n1487), .B0(n1264), .B1(n1475), .Y(n825)
         );
  OAI21XLTS U1098 ( .A0(n826), .A1(n825), .B0(n539), .Y(n824) );
  OAI31X1TS U1099 ( .A0(n826), .A1(n539), .A2(n825), .B0(n824), .Y(
        \mult_x_1/n1090 ) );
  OAI22X1TS U1100 ( .A0(n1646), .A1(n1486), .B0(n1645), .B1(n1494), .Y(n829)
         );
  OAI22X1TS U1101 ( .A0(n1361), .A1(n1488), .B0(n1264), .B1(n1487), .Y(n828)
         );
  OAI21XLTS U1102 ( .A0(n829), .A1(n828), .B0(n539), .Y(n827) );
  OAI31X1TS U1103 ( .A0(n829), .A1(n539), .A2(n828), .B0(n827), .Y(
        \mult_x_1/n1091 ) );
  INVX2TS U1104 ( .A(\mult_x_1/n359 ), .Y(n951) );
  INVX2TS U1105 ( .A(\mult_x_1/n352 ), .Y(n950) );
  INVX2TS U1106 ( .A(n833), .Y(Product[49]) );
  INVX2TS U1107 ( .A(n837), .Y(\mult_x_1/n549 ) );
  XNOR2X1TS U1108 ( .A(n1622), .B(n838), .Y(n839) );
  XOR2XLTS U1109 ( .A(n840), .B(n839), .Y(\mult_x_1/n591 ) );
  INVX2TS U1110 ( .A(n844), .Y(\mult_x_1/n577 ) );
  INVX2TS U1111 ( .A(n848), .Y(\mult_x_1/n563 ) );
  OAI22X1TS U1112 ( .A0(n1554), .A1(n1601), .B0(n1602), .B1(n1553), .Y(n851)
         );
  OAI22X1TS U1113 ( .A0(n927), .A1(n813), .B0(n902), .B1(n1552), .Y(n850) );
  OAI21XLTS U1114 ( .A0(n851), .A1(n850), .B0(n1671), .Y(n849) );
  OAI31X1TS U1115 ( .A0(n851), .A1(n1671), .A2(n850), .B0(n849), .Y(
        \mult_x_1/n1006 ) );
  AOI31XLTS U1116 ( .A0(A[29]), .A1(\mult_x_1/n633 ), .A2(n852), .B0(n1623), 
        .Y(\mult_x_1/n619 ) );
  OAI22X1TS U1117 ( .A0(n723), .A1(n1414), .B0(n727), .B1(n1468), .Y(n855) );
  OAI22X1TS U1118 ( .A0(n1643), .A1(n1435), .B0(n1640), .B1(n1413), .Y(n854)
         );
  OAI21XLTS U1119 ( .A0(n855), .A1(n854), .B0(n1621), .Y(n853) );
  OAI31X1TS U1120 ( .A0(n855), .A1(n1621), .A2(n854), .B0(n853), .Y(
        \mult_x_1/n1034 ) );
  OAI22X1TS U1121 ( .A0(n1186), .A1(n1581), .B0(n1175), .B1(n1580), .Y(n861)
         );
  CLKAND2X2TS U1122 ( .A(n857), .B(n856), .Y(n1188) );
  CLKAND2X2TS U1123 ( .A(n858), .B(n1181), .Y(n1184) );
  OAI22X1TS U1124 ( .A0(n1176), .A1(n1650), .B0(n1177), .B1(n1664), .Y(n860)
         );
  OAI21XLTS U1125 ( .A0(n861), .A1(n860), .B0(n1673), .Y(n859) );
  OAI31X1TS U1126 ( .A0(n861), .A1(n1673), .A2(n860), .B0(n859), .Y(
        \mult_x_1/n1120 ) );
  OAI22X1TS U1127 ( .A0(n989), .A1(n1480), .B0(n1003), .B1(n1479), .Y(n864) );
  OAI22X1TS U1128 ( .A0(n1004), .A1(n1482), .B0(n1005), .B1(n1481), .Y(n863)
         );
  OAI21XLTS U1129 ( .A0(n864), .A1(n863), .B0(n1672), .Y(n862) );
  OAI31X1TS U1130 ( .A0(n864), .A1(n1672), .A2(n863), .B0(n862), .Y(
        \mult_x_1/n1065 ) );
  OAI22X1TS U1131 ( .A0(n989), .A1(n1448), .B0(n1003), .B1(n1482), .Y(n867) );
  OAI22X1TS U1132 ( .A0(n1004), .A1(n1481), .B0(n1005), .B1(n1449), .Y(n866)
         );
  OAI21XLTS U1133 ( .A0(n867), .A1(n866), .B0(n1672), .Y(n865) );
  OAI31X1TS U1134 ( .A0(n867), .A1(n1672), .A2(n866), .B0(n865), .Y(
        \mult_x_1/n1064 ) );
  OAI22X1TS U1135 ( .A0(n989), .A1(n1423), .B0(n1003), .B1(n1481), .Y(n870) );
  OAI22X1TS U1136 ( .A0(n1004), .A1(n1449), .B0(n1005), .B1(n1458), .Y(n869)
         );
  OAI21XLTS U1137 ( .A0(n870), .A1(n869), .B0(n1672), .Y(n868) );
  OAI31X1TS U1138 ( .A0(n870), .A1(n1672), .A2(n869), .B0(n868), .Y(
        \mult_x_1/n1063 ) );
  OAI22X1TS U1139 ( .A0(n723), .A1(n1409), .B0(n727), .B1(n1435), .Y(n873) );
  OAI22X1TS U1140 ( .A0(n1643), .A1(n1413), .B0(n1640), .B1(n1419), .Y(n872)
         );
  OAI21XLTS U1141 ( .A0(n873), .A1(n872), .B0(n1621), .Y(n871) );
  OAI31X1TS U1142 ( .A0(n873), .A1(n1621), .A2(n872), .B0(n871), .Y(
        \mult_x_1/n1035 ) );
  OAI22X1TS U1143 ( .A0(n723), .A1(n1405), .B0(n727), .B1(n1413), .Y(n876) );
  OAI22X1TS U1144 ( .A0(n1643), .A1(n1419), .B0(n1640), .B1(n1501), .Y(n875)
         );
  OAI21XLTS U1145 ( .A0(n876), .A1(n875), .B0(n1621), .Y(n874) );
  OAI31X1TS U1146 ( .A0(n876), .A1(n1621), .A2(n875), .B0(n874), .Y(
        \mult_x_1/n1036 ) );
  OAI22X1TS U1147 ( .A0(n723), .A1(n1418), .B0(n727), .B1(n1419), .Y(n879) );
  OAI22X1TS U1148 ( .A0(n1643), .A1(n1501), .B0(n1640), .B1(n1506), .Y(n878)
         );
  OAI21XLTS U1149 ( .A0(n879), .A1(n878), .B0(n1621), .Y(n877) );
  OAI31X1TS U1150 ( .A0(n879), .A1(n1621), .A2(n878), .B0(n877), .Y(
        \mult_x_1/n1037 ) );
  OAI22X1TS U1151 ( .A0(n723), .A1(n1500), .B0(n727), .B1(n1501), .Y(n882) );
  OAI22X1TS U1152 ( .A0(n1643), .A1(n1506), .B0(n1640), .B1(n1533), .Y(n881)
         );
  OAI21XLTS U1153 ( .A0(n882), .A1(n881), .B0(n1621), .Y(n880) );
  OAI31X1TS U1154 ( .A0(n882), .A1(n1621), .A2(n881), .B0(n880), .Y(
        \mult_x_1/n1038 ) );
  OAI22X1TS U1155 ( .A0(n723), .A1(n1505), .B0(n727), .B1(n1506), .Y(n885) );
  OAI22X1TS U1156 ( .A0(n1643), .A1(n1533), .B0(n1640), .B1(n1552), .Y(n884)
         );
  OAI21XLTS U1157 ( .A0(n885), .A1(n884), .B0(n1621), .Y(n883) );
  OAI31X1TS U1158 ( .A0(n885), .A1(n1621), .A2(n884), .B0(n883), .Y(
        \mult_x_1/n1039 ) );
  OAI22X1TS U1159 ( .A0(n989), .A1(n1444), .B0(n1003), .B1(n1470), .Y(n888) );
  OAI22X1TS U1160 ( .A0(n1004), .A1(n1479), .B0(n1005), .B1(n1482), .Y(n887)
         );
  OAI21XLTS U1161 ( .A0(n888), .A1(n887), .B0(n1672), .Y(n886) );
  OAI31X1TS U1162 ( .A0(n888), .A1(n1672), .A2(n887), .B0(n886), .Y(
        \mult_x_1/n1066 ) );
  OAI22X1TS U1163 ( .A0(n1646), .A1(n1493), .B0(n1645), .B1(n1492), .Y(n891)
         );
  OAI22X1TS U1164 ( .A0(n1361), .A1(n1495), .B0(n1264), .B1(n1494), .Y(n890)
         );
  OAI21XLTS U1165 ( .A0(n891), .A1(n890), .B0(n539), .Y(n889) );
  OAI31X1TS U1166 ( .A0(n891), .A1(n539), .A2(n890), .B0(n889), .Y(
        \mult_x_1/n1093 ) );
  OAI22X1TS U1167 ( .A0(n1646), .A1(n1431), .B0(n1645), .B1(n1495), .Y(n894)
         );
  OAI22X1TS U1168 ( .A0(n1361), .A1(n1494), .B0(n1264), .B1(n1488), .Y(n893)
         );
  OAI21XLTS U1169 ( .A0(n894), .A1(n893), .B0(n539), .Y(n892) );
  OAI31X1TS U1170 ( .A0(n894), .A1(n539), .A2(n893), .B0(n892), .Y(
        \mult_x_1/n1092 ) );
  NOR2XLTS U1171 ( .A(n9), .B(n895), .Y(n1627) );
  OAI222X1TS U1172 ( .A0(n1602), .A1(n1516), .B0(n902), .B1(n23), .C0(n896), 
        .C1(n9), .Y(n1020) );
  AOI21X1TS U1173 ( .A0(A[26]), .A1(n1627), .B0(n1020), .Y(n1030) );
  NAND2X1TS U1174 ( .A(A[26]), .B(n1030), .Y(n901) );
  NOR2XLTS U1175 ( .A(n23), .B(n927), .Y(n898) );
  OAI22X1TS U1176 ( .A0(n9), .A1(n1601), .B0(n1517), .B1(n1602), .Y(n897) );
  AOI211XLTS U1177 ( .A0(n899), .A1(B[2]), .B0(n898), .C0(n897), .Y(n1029) );
  INVX2TS U1178 ( .A(n1029), .Y(n900) );
  NOR2XLTS U1179 ( .A(n901), .B(n900), .Y(\mult_x_1/n645 ) );
  OAI22X1TS U1180 ( .A0(n1527), .A1(n1602), .B0(n23), .B1(n1601), .Y(n905) );
  OAI22X1TS U1181 ( .A0(n1554), .A1(n902), .B0(n29), .B1(n927), .Y(n904) );
  OAI21XLTS U1182 ( .A0(n905), .A1(n904), .B0(n1671), .Y(n903) );
  OAI31X1TS U1183 ( .A0(n905), .A1(n1671), .A2(n904), .B0(n903), .Y(
        \mult_x_1/n1008 ) );
  OAI22X1TS U1184 ( .A0(n989), .A1(n1436), .B0(n1003), .B1(n1435), .Y(n908) );
  OAI22X1TS U1185 ( .A0(n1004), .A1(n1468), .B0(n1005), .B1(n1470), .Y(n907)
         );
  OAI21XLTS U1186 ( .A0(n908), .A1(n907), .B0(n1672), .Y(n906) );
  OAI31X1TS U1187 ( .A0(n908), .A1(n1672), .A2(n907), .B0(n906), .Y(
        \mult_x_1/n1068 ) );
  OAI22X1TS U1188 ( .A0(n989), .A1(n1418), .B0(n1003), .B1(n1506), .Y(n911) );
  OAI22X1TS U1189 ( .A0(n1004), .A1(n1501), .B0(n1005), .B1(n1419), .Y(n910)
         );
  OAI21XLTS U1190 ( .A0(n911), .A1(n910), .B0(n1672), .Y(n909) );
  OAI31X1TS U1191 ( .A0(n911), .A1(n1672), .A2(n910), .B0(n909), .Y(
        \mult_x_1/n1072 ) );
  OAI22X1TS U1192 ( .A0(n989), .A1(n1414), .B0(n1003), .B1(n1413), .Y(n914) );
  OAI22X1TS U1193 ( .A0(n1004), .A1(n1435), .B0(n1005), .B1(n1468), .Y(n913)
         );
  OAI21XLTS U1194 ( .A0(n914), .A1(n913), .B0(n1672), .Y(n912) );
  OAI31X1TS U1195 ( .A0(n914), .A1(n1672), .A2(n913), .B0(n912), .Y(
        \mult_x_1/n1069 ) );
  OAI22X1TS U1196 ( .A0(n989), .A1(n1409), .B0(n1003), .B1(n1419), .Y(n917) );
  OAI22X1TS U1197 ( .A0(n1004), .A1(n1413), .B0(n1005), .B1(n1435), .Y(n916)
         );
  OAI21XLTS U1198 ( .A0(n917), .A1(n916), .B0(n1672), .Y(n915) );
  OAI31X1TS U1199 ( .A0(n917), .A1(n1672), .A2(n916), .B0(n915), .Y(
        \mult_x_1/n1070 ) );
  OAI22X1TS U1200 ( .A0(n989), .A1(n1405), .B0(n1003), .B1(n1501), .Y(n920) );
  OAI22X1TS U1201 ( .A0(n1004), .A1(n1419), .B0(n1005), .B1(n1413), .Y(n919)
         );
  OAI21XLTS U1202 ( .A0(n920), .A1(n919), .B0(n1672), .Y(n918) );
  OAI31X1TS U1203 ( .A0(n920), .A1(n1672), .A2(n919), .B0(n918), .Y(
        \mult_x_1/n1071 ) );
  OAI22X1TS U1204 ( .A0(n989), .A1(n1469), .B0(n1003), .B1(n1468), .Y(n923) );
  OAI22X1TS U1205 ( .A0(n1004), .A1(n1470), .B0(n1005), .B1(n1479), .Y(n922)
         );
  OAI21XLTS U1206 ( .A0(n923), .A1(n922), .B0(n1672), .Y(n921) );
  OAI31X1TS U1207 ( .A0(n923), .A1(n1672), .A2(n922), .B0(n921), .Y(
        \mult_x_1/n1067 ) );
  OAI22X1TS U1208 ( .A0(n989), .A1(n1500), .B0(n1003), .B1(n1533), .Y(n926) );
  OAI22X1TS U1209 ( .A0(n1004), .A1(n1506), .B0(n1005), .B1(n1501), .Y(n925)
         );
  OAI21XLTS U1210 ( .A0(n926), .A1(n925), .B0(n1672), .Y(n924) );
  OAI31X1TS U1211 ( .A0(n926), .A1(n1672), .A2(n925), .B0(n924), .Y(
        \mult_x_1/n1073 ) );
  OAI22X1TS U1212 ( .A0(n29), .A1(n1601), .B0(n1602), .B1(n1537), .Y(n930) );
  OAI22X1TS U1213 ( .A0(n1554), .A1(n927), .B0(n902), .B1(n813), .Y(n929) );
  OAI21XLTS U1214 ( .A0(n930), .A1(n929), .B0(n1671), .Y(n928) );
  OAI31X1TS U1215 ( .A0(n930), .A1(n1671), .A2(n929), .B0(n928), .Y(
        \mult_x_1/n1007 ) );
  OAI22X1TS U1216 ( .A0(n1646), .A1(n1401), .B0(n1645), .B1(n1460), .Y(n933)
         );
  OAI22X1TS U1217 ( .A0(n1361), .A1(n1492), .B0(n1264), .B1(n1495), .Y(n932)
         );
  OAI21XLTS U1218 ( .A0(n933), .A1(n932), .B0(n539), .Y(n931) );
  OAI31X1TS U1219 ( .A0(n933), .A1(n539), .A2(n932), .B0(n931), .Y(
        \mult_x_1/n1094 ) );
  OAI22X1TS U1220 ( .A0(n989), .A1(n1505), .B0(n1003), .B1(n1552), .Y(n936) );
  OAI22X1TS U1221 ( .A0(n1004), .A1(n1533), .B0(n1005), .B1(n1506), .Y(n935)
         );
  OAI21XLTS U1222 ( .A0(n936), .A1(n935), .B0(n1672), .Y(n934) );
  OAI31X1TS U1223 ( .A0(n936), .A1(n1672), .A2(n935), .B0(n934), .Y(
        \mult_x_1/n1074 ) );
  OAI22X1TS U1224 ( .A0(n1186), .A1(n1440), .B0(n1175), .B1(n1454), .Y(n939)
         );
  INVX2TS U1225 ( .A(n1188), .Y(n1176) );
  OAI22X1TS U1226 ( .A0(n1176), .A1(n1560), .B0(n1177), .B1(n1580), .Y(n938)
         );
  OAI21XLTS U1227 ( .A0(n939), .A1(n938), .B0(n1673), .Y(n937) );
  OAI31X1TS U1228 ( .A0(n939), .A1(n1673), .A2(n938), .B0(n937), .Y(
        \mult_x_1/n1122 ) );
  OAI22X1TS U1229 ( .A0(n1186), .A1(n1561), .B0(n1175), .B1(n1560), .Y(n942)
         );
  OAI22X1TS U1230 ( .A0(n1176), .A1(n1580), .B0(n1177), .B1(n1650), .Y(n941)
         );
  OAI21XLTS U1231 ( .A0(n942), .A1(n941), .B0(n1673), .Y(n940) );
  OAI31X1TS U1232 ( .A0(n942), .A1(n1673), .A2(n941), .B0(n940), .Y(
        \mult_x_1/n1121 ) );
  OAI22X1TS U1233 ( .A0(n723), .A1(n1532), .B0(n727), .B1(n1533), .Y(n945) );
  OAI22X1TS U1234 ( .A0(n1643), .A1(n1552), .B0(n1640), .B1(n813), .Y(n944) );
  OAI21XLTS U1235 ( .A0(n945), .A1(n944), .B0(n1621), .Y(n943) );
  OAI31X1TS U1236 ( .A0(n945), .A1(n1621), .A2(n944), .B0(n943), .Y(
        \mult_x_1/n1040 ) );
  OAI22X1TS U1237 ( .A0(n989), .A1(n1532), .B0(n1003), .B1(n813), .Y(n948) );
  OAI22X1TS U1238 ( .A0(n1004), .A1(n1552), .B0(n1005), .B1(n1533), .Y(n947)
         );
  OAI21XLTS U1239 ( .A0(n948), .A1(n947), .B0(n1672), .Y(n946) );
  OAI31X1TS U1240 ( .A0(n948), .A1(n1672), .A2(n947), .B0(n946), .Y(
        \mult_x_1/n1075 ) );
  INVX2TS U1241 ( .A(\mult_x_1/n351 ), .Y(n974) );
  INVX2TS U1242 ( .A(\mult_x_1/n345 ), .Y(n973) );
  INVX2TS U1243 ( .A(n952), .Y(Product[50]) );
  OAI22X1TS U1244 ( .A0(n1186), .A1(n1453), .B0(n1175), .B1(n1475), .Y(n955)
         );
  OAI22X1TS U1245 ( .A0(n1176), .A1(n1454), .B0(n1177), .B1(n1560), .Y(n954)
         );
  OAI21XLTS U1246 ( .A0(n955), .A1(n954), .B0(n1673), .Y(n953) );
  OAI31X1TS U1247 ( .A0(n955), .A1(n1673), .A2(n954), .B0(n953), .Y(
        \mult_x_1/n1123 ) );
  AOI222XLTS U1248 ( .A0(n1182), .A1(n1606), .B0(n1188), .B1(B[31]), .C0(n1), 
        .C1(B[30]), .Y(n956) );
  XOR2XLTS U1249 ( .A(n1673), .B(n956), .Y(\mult_x_1/n1119 ) );
  OAI22X1TS U1250 ( .A0(n1646), .A1(n1459), .B0(n1645), .B1(n1458), .Y(n959)
         );
  OAI22X1TS U1251 ( .A0(n1361), .A1(n1461), .B0(n1264), .B1(n1460), .Y(n958)
         );
  OAI21XLTS U1252 ( .A0(n959), .A1(n958), .B0(n539), .Y(n957) );
  OAI31X1TS U1253 ( .A0(n959), .A1(n539), .A2(n958), .B0(n957), .Y(
        \mult_x_1/n1096 ) );
  OAI22X1TS U1254 ( .A0(n1646), .A1(n1427), .B0(n1645), .B1(n1461), .Y(n962)
         );
  OAI22X1TS U1255 ( .A0(n1361), .A1(n1460), .B0(n1264), .B1(n1492), .Y(n961)
         );
  OAI21XLTS U1256 ( .A0(n962), .A1(n961), .B0(n539), .Y(n960) );
  OAI31X1TS U1257 ( .A0(n962), .A1(n539), .A2(n961), .B0(n960), .Y(
        \mult_x_1/n1095 ) );
  OAI22X1TS U1258 ( .A0(n1554), .A1(n1003), .B0(n989), .B1(n1553), .Y(n965) );
  OAI22X1TS U1259 ( .A0(n1004), .A1(n813), .B0(n1005), .B1(n1552), .Y(n964) );
  OAI21XLTS U1260 ( .A0(n965), .A1(n964), .B0(n1672), .Y(n963) );
  OAI31X1TS U1261 ( .A0(n965), .A1(n1672), .A2(n964), .B0(n963), .Y(
        \mult_x_1/n1076 ) );
  OAI22X1TS U1262 ( .A0(n1186), .A1(n1474), .B0(n1175), .B1(n1488), .Y(n968)
         );
  OAI22X1TS U1263 ( .A0(n1176), .A1(n1487), .B0(n1177), .B1(n1475), .Y(n967)
         );
  OAI21XLTS U1264 ( .A0(n968), .A1(n967), .B0(n1673), .Y(n966) );
  OAI31X1TS U1265 ( .A0(n968), .A1(n1673), .A2(n967), .B0(n966), .Y(
        \mult_x_1/n1125 ) );
  OAI22X1TS U1266 ( .A0(n1186), .A1(n1397), .B0(n1175), .B1(n1487), .Y(n971)
         );
  OAI22X1TS U1267 ( .A0(n1176), .A1(n1475), .B0(n1177), .B1(n1454), .Y(n970)
         );
  OAI21XLTS U1268 ( .A0(n971), .A1(n970), .B0(n1673), .Y(n969) );
  OAI31X1TS U1269 ( .A0(n971), .A1(n1673), .A2(n970), .B0(n969), .Y(
        \mult_x_1/n1124 ) );
  INVX2TS U1270 ( .A(\mult_x_1/n344 ), .Y(n995) );
  INVX2TS U1271 ( .A(\mult_x_1/n337 ), .Y(n994) );
  INVX2TS U1272 ( .A(n975), .Y(Product[51]) );
  OAI22X1TS U1273 ( .A0(n1646), .A1(n1393), .B0(n1645), .B1(n1449), .Y(n978)
         );
  OAI22X1TS U1274 ( .A0(n1361), .A1(n1458), .B0(n1264), .B1(n1461), .Y(n977)
         );
  OAI21XLTS U1275 ( .A0(n978), .A1(n977), .B0(n539), .Y(n976) );
  OAI31X1TS U1276 ( .A0(n978), .A1(n539), .A2(n977), .B0(n976), .Y(
        \mult_x_1/n1097 ) );
  OAI22X1TS U1277 ( .A0(n29), .A1(n1003), .B0(n989), .B1(n1537), .Y(n981) );
  OAI22X1TS U1278 ( .A0(n1554), .A1(n1004), .B0(n1005), .B1(n813), .Y(n980) );
  OAI21XLTS U1279 ( .A0(n981), .A1(n980), .B0(n1672), .Y(n979) );
  OAI31X1TS U1280 ( .A0(n981), .A1(n1672), .A2(n980), .B0(n979), .Y(
        \mult_x_1/n1077 ) );
  OAI22X1TS U1281 ( .A0(n1186), .A1(n1486), .B0(n1175), .B1(n1494), .Y(n984)
         );
  OAI22X1TS U1282 ( .A0(n1176), .A1(n1488), .B0(n1177), .B1(n1487), .Y(n983)
         );
  OAI21XLTS U1283 ( .A0(n984), .A1(n983), .B0(n1673), .Y(n982) );
  OAI31X1TS U1284 ( .A0(n984), .A1(n1673), .A2(n983), .B0(n982), .Y(
        \mult_x_1/n1126 ) );
  NAND2X1TS U1285 ( .A(B[0]), .B(n985), .Y(n1351) );
  AOI222XLTS U1286 ( .A0(B[1]), .A1(n987), .B0(B[0]), .B1(n991), .C0(n1183), 
        .C1(n540), .Y(n1352) );
  OAI21XLTS U1287 ( .A0(n1672), .A1(n1351), .B0(n1352), .Y(n1354) );
  AOI22X1TS U1288 ( .A0(B[2]), .A1(n987), .B0(B[0]), .B1(n986), .Y(n988) );
  OAI21XLTS U1289 ( .A0(n1517), .A1(n989), .B0(n988), .Y(n990) );
  AOI21X1TS U1290 ( .A0(B[1]), .A1(n991), .B0(n990), .Y(n1356) );
  NAND2X1TS U1291 ( .A(A[20]), .B(n1356), .Y(n992) );
  NOR2XLTS U1292 ( .A(n1354), .B(n992), .Y(\mult_x_1/n714 ) );
  INVX2TS U1293 ( .A(\mult_x_1/n336 ), .Y(n1070) );
  INVX2TS U1294 ( .A(\mult_x_1/n332 ), .Y(n1069) );
  INVX2TS U1295 ( .A(n996), .Y(Product[52]) );
  AOI2BB2XLTS U1296 ( .B0(A[11]), .B1(A[10]), .A0N(A[10]), .A1N(A[11]), .Y(
        n999) );
  OAI2BB2XLTS U1297 ( .B0(n1674), .B1(A[9]), .A0N(A[9]), .A1N(n1674), .Y(n997)
         );
  NAND2X1TS U1298 ( .A(n999), .B(n997), .Y(n1164) );
  CLKBUFX2TS U1299 ( .A(n1164), .Y(n1654) );
  OAI22X1TS U1300 ( .A0(n1654), .A1(n1581), .B0(n1518), .B1(n1664), .Y(n1002)
         );
  XNOR2X1TS U1301 ( .A(A[10]), .B(A[9]), .Y(n998) );
  INVX2TS U1302 ( .A(n997), .Y(n1515) );
  NAND3XLTS U1303 ( .A(n999), .B(n1515), .C(n998), .Y(n1651) );
  CLKBUFX2TS U1304 ( .A(n1651), .Y(n1648) );
  OAI22X1TS U1305 ( .A0(n1652), .A1(n1650), .B0(n1648), .B1(n1580), .Y(n1001)
         );
  OAI21XLTS U1306 ( .A0(n1002), .A1(n1001), .B0(n1638), .Y(n1000) );
  OAI31X1TS U1307 ( .A0(n1002), .A1(n1638), .A2(n1001), .B0(n1000), .Y(
        \mult_x_1/n1155 ) );
  OAI22X1TS U1308 ( .A0(n1527), .A1(n989), .B0(n23), .B1(n1003), .Y(n1008) );
  OAI22X1TS U1309 ( .A0(n1554), .A1(n1005), .B0(n29), .B1(n1004), .Y(n1007) );
  OAI21XLTS U1310 ( .A0(n1008), .A1(n1007), .B0(n1672), .Y(n1006) );
  OAI31X1TS U1311 ( .A0(n1008), .A1(n1672), .A2(n1007), .B0(n1006), .Y(
        \mult_x_1/n1078 ) );
  OAI22X1TS U1312 ( .A0(n723), .A1(n1537), .B0(n727), .B1(n813), .Y(n1011) );
  OAI22X1TS U1313 ( .A0(n1554), .A1(n1643), .B0(n29), .B1(n1640), .Y(n1010) );
  OAI21XLTS U1314 ( .A0(n1011), .A1(n1010), .B0(A[23]), .Y(n1009) );
  OAI31X1TS U1315 ( .A0(n1011), .A1(A[23]), .A2(n1010), .B0(n1009), .Y(n1033)
         );
  NOR2XLTS U1316 ( .A(n9), .B(n1012), .Y(\mult_x_1/n705 ) );
  OAI222X1TS U1317 ( .A0(n723), .A1(n1516), .B0(n727), .B1(n23), .C0(n1643), 
        .C1(n9), .Y(n1610) );
  AOI21X1TS U1318 ( .A0(A[23]), .A1(\mult_x_1/n705 ), .B0(n1610), .Y(n1609) );
  NAND2X1TS U1319 ( .A(A[23]), .B(n1609), .Y(n1016) );
  OAI22X1TS U1320 ( .A0(n29), .A1(n727), .B0(n1517), .B1(n723), .Y(n1014) );
  OAI22X1TS U1321 ( .A0(n23), .A1(n1643), .B0(n9), .B1(n1640), .Y(n1013) );
  NOR2XLTS U1322 ( .A(n1014), .B(n1013), .Y(n1027) );
  INVX2TS U1323 ( .A(n1027), .Y(n1015) );
  NOR2XLTS U1324 ( .A(n1016), .B(n1015), .Y(n1628) );
  OAI22X1TS U1325 ( .A0(n1554), .A1(n727), .B0(n1527), .B1(n723), .Y(n1019) );
  OAI22X1TS U1326 ( .A0(n29), .A1(n1643), .B0(n23), .B1(n1640), .Y(n1018) );
  OAI21XLTS U1327 ( .A0(n1019), .A1(n1018), .B0(n1621), .Y(n1017) );
  OAI31X1TS U1328 ( .A0(n1019), .A1(n1621), .A2(n1018), .B0(n1017), .Y(n1630)
         );
  OAI21XLTS U1329 ( .A0(n1628), .A1(n1627), .B0(n1630), .Y(n1032) );
  NOR2BX1TS U1330 ( .AN(n1627), .B(n1671), .Y(n1021) );
  AO21XLTS U1331 ( .A0(n1021), .A1(n1020), .B0(n1030), .Y(n1031) );
  INVX2TS U1332 ( .A(n1022), .Y(\mult_x_1/n657 ) );
  OAI22X1TS U1333 ( .A0(n1646), .A1(n1423), .B0(n1645), .B1(n1481), .Y(n1025)
         );
  OAI22X1TS U1334 ( .A0(n1361), .A1(n1449), .B0(n1264), .B1(n1458), .Y(n1024)
         );
  OAI21XLTS U1335 ( .A0(n1025), .A1(n1024), .B0(n539), .Y(n1023) );
  OAI31X1TS U1336 ( .A0(n1025), .A1(n539), .A2(n1024), .B0(n1023), .Y(
        \mult_x_1/n1098 ) );
  NOR3XLTS U1337 ( .A(n1027), .B(n1609), .C(n1621), .Y(n1026) );
  AOI211XLTS U1338 ( .A0(n1027), .A1(n1621), .B0(n1628), .C0(n1026), .Y(
        \mult_x_1/n683 ) );
  OAI21XLTS U1339 ( .A0(n1030), .A1(n1671), .B0(n1029), .Y(n1028) );
  OAI31X1TS U1340 ( .A0(n1030), .A1(n1029), .A2(n1671), .B0(n1028), .Y(n1086)
         );
  OAI22X1TS U1341 ( .A0(n723), .A1(n1553), .B0(n727), .B1(n1552), .Y(n1036) );
  OAI22X1TS U1342 ( .A0(n1554), .A1(n1640), .B0(n1643), .B1(n813), .Y(n1035)
         );
  OAI21XLTS U1343 ( .A0(n1036), .A1(n1035), .B0(A[23]), .Y(n1034) );
  OAI31X1TS U1344 ( .A0(n1036), .A1(A[23]), .A2(n1035), .B0(n1034), .Y(n1084)
         );
  INVX2TS U1345 ( .A(n1037), .Y(\mult_x_1/n643 ) );
  OAI22X1TS U1346 ( .A0(n1646), .A1(n1444), .B0(n1645), .B1(n1470), .Y(n1040)
         );
  OAI22X1TS U1347 ( .A0(n1346), .A1(n1479), .B0(n1264), .B1(n1482), .Y(n1039)
         );
  OAI21XLTS U1348 ( .A0(n1040), .A1(n1039), .B0(n539), .Y(n1038) );
  OAI31X1TS U1349 ( .A0(n1040), .A1(n539), .A2(n1039), .B0(n1038), .Y(
        \mult_x_1/n1101 ) );
  OAI22X1TS U1350 ( .A0(n1646), .A1(n1418), .B0(n1645), .B1(n1506), .Y(n1043)
         );
  OAI22X1TS U1351 ( .A0(n1346), .A1(n1501), .B0(n1264), .B1(n1419), .Y(n1042)
         );
  OAI21XLTS U1352 ( .A0(n1043), .A1(n1042), .B0(n539), .Y(n1041) );
  OAI31X1TS U1353 ( .A0(n1043), .A1(n539), .A2(n1042), .B0(n1041), .Y(
        \mult_x_1/n1107 ) );
  OAI22X1TS U1354 ( .A0(n1646), .A1(n1414), .B0(n1645), .B1(n1413), .Y(n1046)
         );
  OAI22X1TS U1355 ( .A0(n1346), .A1(n1435), .B0(n1264), .B1(n1468), .Y(n1045)
         );
  OAI21XLTS U1356 ( .A0(n1046), .A1(n1045), .B0(n539), .Y(n1044) );
  OAI31X1TS U1357 ( .A0(n1046), .A1(n539), .A2(n1045), .B0(n1044), .Y(
        \mult_x_1/n1104 ) );
  OAI22X1TS U1358 ( .A0(n1646), .A1(n1405), .B0(n1645), .B1(n1501), .Y(n1049)
         );
  OAI22X1TS U1359 ( .A0(n1346), .A1(n1419), .B0(n1264), .B1(n1413), .Y(n1048)
         );
  OAI21XLTS U1360 ( .A0(n1049), .A1(n1048), .B0(n539), .Y(n1047) );
  OAI31X1TS U1361 ( .A0(n1049), .A1(n539), .A2(n1048), .B0(n1047), .Y(
        \mult_x_1/n1106 ) );
  OAI22X1TS U1362 ( .A0(n1646), .A1(n1469), .B0(n1645), .B1(n1468), .Y(n1052)
         );
  OAI22X1TS U1363 ( .A0(n1346), .A1(n1470), .B0(n1264), .B1(n1479), .Y(n1051)
         );
  OAI21XLTS U1364 ( .A0(n1052), .A1(n1051), .B0(n539), .Y(n1050) );
  OAI31X1TS U1365 ( .A0(n1052), .A1(n539), .A2(n1051), .B0(n1050), .Y(
        \mult_x_1/n1102 ) );
  OAI22X1TS U1366 ( .A0(n1646), .A1(n1436), .B0(n1645), .B1(n1435), .Y(n1055)
         );
  OAI22X1TS U1367 ( .A0(n1346), .A1(n1468), .B0(n1264), .B1(n1470), .Y(n1054)
         );
  OAI21XLTS U1368 ( .A0(n1055), .A1(n1054), .B0(n539), .Y(n1053) );
  OAI31X1TS U1369 ( .A0(n1055), .A1(n539), .A2(n1054), .B0(n1053), .Y(
        \mult_x_1/n1103 ) );
  OAI22X1TS U1370 ( .A0(n1646), .A1(n1448), .B0(n1645), .B1(n1482), .Y(n1058)
         );
  OAI22X1TS U1371 ( .A0(n1346), .A1(n1481), .B0(n1264), .B1(n1449), .Y(n1057)
         );
  OAI21XLTS U1372 ( .A0(n1058), .A1(n1057), .B0(n539), .Y(n1056) );
  OAI31X1TS U1373 ( .A0(n1058), .A1(n539), .A2(n1057), .B0(n1056), .Y(
        \mult_x_1/n1099 ) );
  OAI22X1TS U1374 ( .A0(n1646), .A1(n1480), .B0(n1645), .B1(n1479), .Y(n1061)
         );
  OAI22X1TS U1375 ( .A0(n1346), .A1(n1482), .B0(n1264), .B1(n1481), .Y(n1060)
         );
  OAI21XLTS U1376 ( .A0(n1061), .A1(n1060), .B0(n539), .Y(n1059) );
  OAI31X1TS U1377 ( .A0(n1061), .A1(n539), .A2(n1060), .B0(n1059), .Y(
        \mult_x_1/n1100 ) );
  OAI22X1TS U1378 ( .A0(n1646), .A1(n1409), .B0(n1645), .B1(n1419), .Y(n1064)
         );
  OAI22X1TS U1379 ( .A0(n1346), .A1(n1413), .B0(n1264), .B1(n1435), .Y(n1063)
         );
  OAI21XLTS U1380 ( .A0(n1064), .A1(n1063), .B0(n539), .Y(n1062) );
  OAI31X1TS U1381 ( .A0(n1064), .A1(n539), .A2(n1063), .B0(n1062), .Y(
        \mult_x_1/n1105 ) );
  OAI22X1TS U1382 ( .A0(n1646), .A1(n1500), .B0(n1645), .B1(n1533), .Y(n1067)
         );
  OAI22X1TS U1383 ( .A0(n1346), .A1(n1506), .B0(n1264), .B1(n1501), .Y(n1066)
         );
  OAI21XLTS U1384 ( .A0(n1067), .A1(n1066), .B0(n539), .Y(n1065) );
  OAI31X1TS U1385 ( .A0(n1067), .A1(n539), .A2(n1066), .B0(n1065), .Y(
        \mult_x_1/n1108 ) );
  INVX2TS U1386 ( .A(\mult_x_1/n331 ), .Y(n1159) );
  INVX2TS U1387 ( .A(\mult_x_1/n326 ), .Y(n1158) );
  INVX2TS U1388 ( .A(n1071), .Y(Product[53]) );
  OAI22X1TS U1389 ( .A0(n1186), .A1(n1493), .B0(n1175), .B1(n1492), .Y(n1074)
         );
  OAI22X1TS U1390 ( .A0(n1176), .A1(n1495), .B0(n1177), .B1(n1494), .Y(n1073)
         );
  OAI21XLTS U1391 ( .A0(n1074), .A1(n1073), .B0(n1673), .Y(n1072) );
  OAI31X1TS U1392 ( .A0(n1074), .A1(n1673), .A2(n1073), .B0(n1072), .Y(
        \mult_x_1/n1128 ) );
  OAI22X1TS U1393 ( .A0(n1186), .A1(n1401), .B0(n1175), .B1(n1460), .Y(n1077)
         );
  OAI22X1TS U1394 ( .A0(n1176), .A1(n1492), .B0(n1177), .B1(n1495), .Y(n1076)
         );
  OAI21XLTS U1395 ( .A0(n1077), .A1(n1076), .B0(n1673), .Y(n1075) );
  OAI31X1TS U1396 ( .A0(n1077), .A1(n1673), .A2(n1076), .B0(n1075), .Y(
        \mult_x_1/n1129 ) );
  OAI22X1TS U1397 ( .A0(n1186), .A1(n1431), .B0(n1175), .B1(n1495), .Y(n1080)
         );
  OAI22X1TS U1398 ( .A0(n1176), .A1(n1494), .B0(n1177), .B1(n1488), .Y(n1079)
         );
  OAI21XLTS U1399 ( .A0(n1080), .A1(n1079), .B0(n1673), .Y(n1078) );
  OAI31X1TS U1400 ( .A0(n1080), .A1(n1673), .A2(n1079), .B0(n1078), .Y(
        \mult_x_1/n1127 ) );
  OAI22X1TS U1401 ( .A0(n1646), .A1(n1505), .B0(n1645), .B1(n1552), .Y(n1083)
         );
  OAI22X1TS U1402 ( .A0(n1346), .A1(n1533), .B0(n1264), .B1(n1506), .Y(n1082)
         );
  OAI21XLTS U1403 ( .A0(n1083), .A1(n1082), .B0(n539), .Y(n1081) );
  OAI31X1TS U1404 ( .A0(n1083), .A1(n539), .A2(n1082), .B0(n1081), .Y(
        \mult_x_1/n1109 ) );
  INVX2TS U1405 ( .A(n1087), .Y(\mult_x_1/n644 ) );
  OAI22X1TS U1406 ( .A0(n1186), .A1(n1427), .B0(n1175), .B1(n1461), .Y(n1090)
         );
  OAI22X1TS U1407 ( .A0(n1176), .A1(n1460), .B0(n1177), .B1(n1492), .Y(n1089)
         );
  OAI21XLTS U1408 ( .A0(n1090), .A1(n1089), .B0(n1673), .Y(n1088) );
  OAI31X1TS U1409 ( .A0(n1090), .A1(n1673), .A2(n1089), .B0(n1088), .Y(
        \mult_x_1/n1130 ) );
  OAI22X1TS U1410 ( .A0(n1186), .A1(n1459), .B0(n1175), .B1(n1458), .Y(n1093)
         );
  OAI22X1TS U1411 ( .A0(n1176), .A1(n1461), .B0(n1177), .B1(n1460), .Y(n1092)
         );
  OAI21XLTS U1412 ( .A0(n1093), .A1(n1092), .B0(n1673), .Y(n1091) );
  OAI31X1TS U1413 ( .A0(n1093), .A1(n1673), .A2(n1092), .B0(n1091), .Y(
        \mult_x_1/n1131 ) );
  OAI22X1TS U1414 ( .A0(n1186), .A1(n1393), .B0(n1175), .B1(n1449), .Y(n1096)
         );
  INVX2TS U1415 ( .A(n1184), .Y(n1177) );
  OAI22X1TS U1416 ( .A0(n1176), .A1(n1458), .B0(n1177), .B1(n1461), .Y(n1095)
         );
  OAI21XLTS U1417 ( .A0(n1096), .A1(n1095), .B0(n1673), .Y(n1094) );
  OAI31X1TS U1418 ( .A0(n1096), .A1(n1673), .A2(n1095), .B0(n1094), .Y(
        \mult_x_1/n1132 ) );
  OAI22X1TS U1419 ( .A0(n1186), .A1(n1448), .B0(n1175), .B1(n1482), .Y(n1099)
         );
  OAI22X1TS U1420 ( .A0(n1176), .A1(n1481), .B0(n1177), .B1(n1449), .Y(n1098)
         );
  OAI21XLTS U1421 ( .A0(n1099), .A1(n1098), .B0(n1673), .Y(n1097) );
  OAI31X1TS U1422 ( .A0(n1099), .A1(n1673), .A2(n1098), .B0(n1097), .Y(
        \mult_x_1/n1134 ) );
  OAI22X1TS U1423 ( .A0(n1186), .A1(n1480), .B0(n1175), .B1(n1479), .Y(n1102)
         );
  OAI22X1TS U1424 ( .A0(n1176), .A1(n1482), .B0(n1177), .B1(n1481), .Y(n1101)
         );
  OAI21XLTS U1425 ( .A0(n1102), .A1(n1101), .B0(n1673), .Y(n1100) );
  OAI31X1TS U1426 ( .A0(n1102), .A1(n1673), .A2(n1101), .B0(n1100), .Y(
        \mult_x_1/n1135 ) );
  OAI22X1TS U1427 ( .A0(n1186), .A1(n1405), .B0(n1175), .B1(n1501), .Y(n1105)
         );
  OAI22X1TS U1428 ( .A0(n1176), .A1(n1419), .B0(n1177), .B1(n1413), .Y(n1104)
         );
  OAI21XLTS U1429 ( .A0(n1105), .A1(n1104), .B0(n1673), .Y(n1103) );
  OAI31X1TS U1430 ( .A0(n1105), .A1(n1673), .A2(n1104), .B0(n1103), .Y(
        \mult_x_1/n1141 ) );
  OAI22X1TS U1431 ( .A0(n1186), .A1(n1436), .B0(n1175), .B1(n1435), .Y(n1108)
         );
  OAI22X1TS U1432 ( .A0(n1176), .A1(n1468), .B0(n1177), .B1(n1470), .Y(n1107)
         );
  OAI21XLTS U1433 ( .A0(n1108), .A1(n1107), .B0(n1673), .Y(n1106) );
  OAI31X1TS U1434 ( .A0(n1108), .A1(n1673), .A2(n1107), .B0(n1106), .Y(
        \mult_x_1/n1138 ) );
  OAI22X1TS U1435 ( .A0(n1186), .A1(n1423), .B0(n1175), .B1(n1481), .Y(n1111)
         );
  OAI22X1TS U1436 ( .A0(n1176), .A1(n1449), .B0(n1177), .B1(n1458), .Y(n1110)
         );
  OAI21XLTS U1437 ( .A0(n1111), .A1(n1110), .B0(n1673), .Y(n1109) );
  OAI31X1TS U1438 ( .A0(n1111), .A1(n1673), .A2(n1110), .B0(n1109), .Y(
        \mult_x_1/n1133 ) );
  OAI22X1TS U1439 ( .A0(n1186), .A1(n1414), .B0(n1175), .B1(n1413), .Y(n1114)
         );
  OAI22X1TS U1440 ( .A0(n1176), .A1(n1435), .B0(n1177), .B1(n1468), .Y(n1113)
         );
  OAI21XLTS U1441 ( .A0(n1114), .A1(n1113), .B0(n1673), .Y(n1112) );
  OAI31X1TS U1442 ( .A0(n1114), .A1(n1673), .A2(n1113), .B0(n1112), .Y(
        \mult_x_1/n1139 ) );
  OAI22X1TS U1443 ( .A0(n1186), .A1(n1409), .B0(n1175), .B1(n1419), .Y(n1117)
         );
  OAI22X1TS U1444 ( .A0(n1176), .A1(n1413), .B0(n1177), .B1(n1435), .Y(n1116)
         );
  OAI21XLTS U1445 ( .A0(n1117), .A1(n1116), .B0(n1673), .Y(n1115) );
  OAI31X1TS U1446 ( .A0(n1117), .A1(n1673), .A2(n1116), .B0(n1115), .Y(
        \mult_x_1/n1140 ) );
  OAI22X1TS U1447 ( .A0(n1186), .A1(n1444), .B0(n1175), .B1(n1470), .Y(n1120)
         );
  OAI22X1TS U1448 ( .A0(n1176), .A1(n1479), .B0(n1177), .B1(n1482), .Y(n1119)
         );
  OAI21XLTS U1449 ( .A0(n1120), .A1(n1119), .B0(n1673), .Y(n1118) );
  OAI31X1TS U1450 ( .A0(n1120), .A1(n1673), .A2(n1119), .B0(n1118), .Y(
        \mult_x_1/n1136 ) );
  OAI22X1TS U1451 ( .A0(n1186), .A1(n1469), .B0(n1175), .B1(n1468), .Y(n1123)
         );
  OAI22X1TS U1452 ( .A0(n1176), .A1(n1470), .B0(n1177), .B1(n1479), .Y(n1122)
         );
  OAI21XLTS U1453 ( .A0(n1123), .A1(n1122), .B0(n1673), .Y(n1121) );
  OAI31X1TS U1454 ( .A0(n1123), .A1(n1673), .A2(n1122), .B0(n1121), .Y(
        \mult_x_1/n1137 ) );
  OAI22X1TS U1455 ( .A0(n1186), .A1(n1418), .B0(n1175), .B1(n1506), .Y(n1126)
         );
  OAI22X1TS U1456 ( .A0(n1176), .A1(n1501), .B0(n1177), .B1(n1419), .Y(n1125)
         );
  OAI21XLTS U1457 ( .A0(n1126), .A1(n1125), .B0(n1673), .Y(n1124) );
  OAI31X1TS U1458 ( .A0(n1126), .A1(n1673), .A2(n1125), .B0(n1124), .Y(
        \mult_x_1/n1142 ) );
  OAI22X1TS U1459 ( .A0(n1186), .A1(n1500), .B0(n1175), .B1(n1533), .Y(n1129)
         );
  OAI22X1TS U1460 ( .A0(n1176), .A1(n1506), .B0(n1177), .B1(n1501), .Y(n1128)
         );
  OAI21XLTS U1461 ( .A0(n1129), .A1(n1128), .B0(n1673), .Y(n1127) );
  OAI31X1TS U1462 ( .A0(n1129), .A1(n1673), .A2(n1128), .B0(n1127), .Y(
        \mult_x_1/n1143 ) );
  OAI22X1TS U1463 ( .A0(n1164), .A1(n1561), .B0(n1518), .B1(n1650), .Y(n1132)
         );
  OAI22X1TS U1464 ( .A0(n1652), .A1(n1580), .B0(n1651), .B1(n1560), .Y(n1131)
         );
  OAI21XLTS U1465 ( .A0(n1132), .A1(n1131), .B0(n1638), .Y(n1130) );
  OAI31X1TS U1466 ( .A0(n1132), .A1(n1638), .A2(n1131), .B0(n1130), .Y(
        \mult_x_1/n1156 ) );
  OAI22X1TS U1467 ( .A0(n1164), .A1(n1440), .B0(n1518), .B1(n1580), .Y(n1135)
         );
  OAI22X1TS U1468 ( .A0(n1652), .A1(n1560), .B0(n1651), .B1(n1454), .Y(n1134)
         );
  OAI21XLTS U1469 ( .A0(n1135), .A1(n1134), .B0(n1638), .Y(n1133) );
  OAI31X1TS U1470 ( .A0(n1135), .A1(n1638), .A2(n1134), .B0(n1133), .Y(
        \mult_x_1/n1157 ) );
  OAI22X1TS U1471 ( .A0(n1646), .A1(n1532), .B0(n1645), .B1(n813), .Y(n1138)
         );
  OAI22X1TS U1472 ( .A0(n1361), .A1(n1552), .B0(n1264), .B1(n1533), .Y(n1137)
         );
  OAI21XLTS U1473 ( .A0(n1138), .A1(n1137), .B0(n539), .Y(n1136) );
  OAI31X1TS U1474 ( .A0(n1138), .A1(n539), .A2(n1137), .B0(n1136), .Y(
        \mult_x_1/n1110 ) );
  OAI22X1TS U1475 ( .A0(n1186), .A1(n1505), .B0(n1175), .B1(n1552), .Y(n1141)
         );
  OAI22X1TS U1476 ( .A0(n1176), .A1(n1533), .B0(n1177), .B1(n1506), .Y(n1140)
         );
  OAI21XLTS U1477 ( .A0(n1141), .A1(n1140), .B0(n1673), .Y(n1139) );
  OAI31X1TS U1478 ( .A0(n1141), .A1(n1673), .A2(n1140), .B0(n1139), .Y(
        \mult_x_1/n1144 ) );
  OAI22X1TS U1479 ( .A0(n1164), .A1(n1453), .B0(n1518), .B1(n1560), .Y(n1144)
         );
  OAI22X1TS U1480 ( .A0(n1652), .A1(n1454), .B0(n1651), .B1(n1475), .Y(n1143)
         );
  OAI21XLTS U1481 ( .A0(n1144), .A1(n1143), .B0(n1638), .Y(n1142) );
  OAI31X1TS U1482 ( .A0(n1144), .A1(n1638), .A2(n1143), .B0(n1142), .Y(
        \mult_x_1/n1158 ) );
  OAI22X1TS U1483 ( .A0(n1186), .A1(n1532), .B0(n1175), .B1(n813), .Y(n1147)
         );
  OAI22X1TS U1484 ( .A0(n1176), .A1(n1552), .B0(n1177), .B1(n1533), .Y(n1146)
         );
  OAI21XLTS U1485 ( .A0(n1147), .A1(n1146), .B0(n1673), .Y(n1145) );
  OAI31X1TS U1486 ( .A0(n1147), .A1(n1673), .A2(n1146), .B0(n1145), .Y(
        \mult_x_1/n1145 ) );
  OAI22X1TS U1487 ( .A0(n1164), .A1(n1397), .B0(n1518), .B1(n1454), .Y(n1150)
         );
  OAI22X1TS U1488 ( .A0(n1652), .A1(n1475), .B0(n1651), .B1(n1487), .Y(n1149)
         );
  OAI21XLTS U1489 ( .A0(n1150), .A1(n1149), .B0(n1638), .Y(n1148) );
  OAI31X1TS U1490 ( .A0(n1150), .A1(n1638), .A2(n1149), .B0(n1148), .Y(
        \mult_x_1/n1159 ) );
  OAI22X1TS U1491 ( .A0(n1164), .A1(n1474), .B0(n1518), .B1(n1475), .Y(n1153)
         );
  OAI22X1TS U1492 ( .A0(n1652), .A1(n1487), .B0(n1651), .B1(n1488), .Y(n1152)
         );
  OAI21XLTS U1493 ( .A0(n1153), .A1(n1152), .B0(n1638), .Y(n1151) );
  OAI31X1TS U1494 ( .A0(n1153), .A1(n1638), .A2(n1152), .B0(n1151), .Y(
        \mult_x_1/n1160 ) );
  OAI22X1TS U1495 ( .A0(n1554), .A1(n1175), .B0(n1186), .B1(n1553), .Y(n1156)
         );
  OAI22X1TS U1496 ( .A0(n1176), .A1(n813), .B0(n1177), .B1(n1552), .Y(n1155)
         );
  OAI21XLTS U1497 ( .A0(n1156), .A1(n1155), .B0(n1673), .Y(n1154) );
  OAI31X1TS U1498 ( .A0(n1156), .A1(n1673), .A2(n1155), .B0(n1154), .Y(
        \mult_x_1/n1146 ) );
  INVX2TS U1499 ( .A(\mult_x_1/n325 ), .Y(n1170) );
  INVX2TS U1500 ( .A(\mult_x_1/n319 ), .Y(n1169) );
  INVX2TS U1501 ( .A(n1160), .Y(Product[54]) );
  OAI22X1TS U1502 ( .A0(n29), .A1(n1175), .B0(n1186), .B1(n1537), .Y(n1163) );
  OAI22X1TS U1503 ( .A0(n1554), .A1(n1176), .B0(n1177), .B1(n813), .Y(n1162)
         );
  OAI21XLTS U1504 ( .A0(n1163), .A1(n1162), .B0(n1673), .Y(n1161) );
  OAI31X1TS U1505 ( .A0(n1163), .A1(n1673), .A2(n1162), .B0(n1161), .Y(
        \mult_x_1/n1147 ) );
  OAI22X1TS U1506 ( .A0(n1164), .A1(n1486), .B0(n1518), .B1(n1487), .Y(n1167)
         );
  OAI22X1TS U1507 ( .A0(n1652), .A1(n1488), .B0(n1648), .B1(n1494), .Y(n1166)
         );
  OAI21XLTS U1508 ( .A0(n1167), .A1(n1166), .B0(n1638), .Y(n1165) );
  OAI31X1TS U1509 ( .A0(n1167), .A1(n1638), .A2(n1166), .B0(n1165), .Y(
        \mult_x_1/n1161 ) );
  INVX2TS U1510 ( .A(\mult_x_1/n318 ), .Y(n1258) );
  INVX2TS U1511 ( .A(\mult_x_1/n315 ), .Y(n1257) );
  INVX2TS U1512 ( .A(n1171), .Y(Product[55]) );
  OAI22X1TS U1513 ( .A0(n1657), .A1(n1581), .B0(n1656), .B1(n1580), .Y(n1174)
         );
  OAI22X1TS U1514 ( .A0(n1528), .A1(n1650), .B0(n1279), .B1(n1664), .Y(n1173)
         );
  OAI21XLTS U1515 ( .A0(n1174), .A1(n1173), .B0(n1674), .Y(n1172) );
  OAI31X1TS U1516 ( .A0(n1174), .A1(n1674), .A2(n1173), .B0(n1172), .Y(
        \mult_x_1/n1190 ) );
  OAI22X1TS U1517 ( .A0(n1527), .A1(n1186), .B0(n23), .B1(n1175), .Y(n1180) );
  OAI22X1TS U1518 ( .A0(n1554), .A1(n1177), .B0(n29), .B1(n1176), .Y(n1179) );
  OAI21XLTS U1519 ( .A0(n1180), .A1(n1179), .B0(n1673), .Y(n1178) );
  OAI31X1TS U1520 ( .A0(n1180), .A1(n1673), .A2(n1179), .B0(n1178), .Y(
        \mult_x_1/n1148 ) );
  NAND2X1TS U1521 ( .A(B[0]), .B(n1181), .Y(n1542) );
  AOI222XLTS U1522 ( .A0(B[1]), .A1(n1184), .B0(B[0]), .B1(n1188), .C0(n1183), 
        .C1(n1182), .Y(n1543) );
  OAI21XLTS U1523 ( .A0(n1673), .A1(n1542), .B0(n1543), .Y(n1545) );
  AOI22X1TS U1524 ( .A0(B[2]), .A1(n1184), .B0(B[0]), .B1(n1), .Y(n1185) );
  OAI21XLTS U1525 ( .A0(n1517), .A1(n1186), .B0(n1185), .Y(n1187) );
  AOI21X1TS U1526 ( .A0(B[1]), .A1(n1188), .B0(n1187), .Y(n1547) );
  NAND2X1TS U1527 ( .A(A[14]), .B(n1547), .Y(n1189) );
  NOR2XLTS U1528 ( .A(n1545), .B(n1189), .Y(\mult_x_1/n765 ) );
  OAI22X1TS U1529 ( .A0(n1654), .A1(n1431), .B0(n1518), .B1(n1488), .Y(n1192)
         );
  OAI22X1TS U1530 ( .A0(n1652), .A1(n1494), .B0(n1648), .B1(n1495), .Y(n1191)
         );
  OAI21XLTS U1531 ( .A0(n1192), .A1(n1191), .B0(n1638), .Y(n1190) );
  OAI31X1TS U1532 ( .A0(n1192), .A1(n1638), .A2(n1191), .B0(n1190), .Y(
        \mult_x_1/n1162 ) );
  OAI22X1TS U1533 ( .A0(n1654), .A1(n1405), .B0(n1518), .B1(n1413), .Y(n1195)
         );
  OAI22X1TS U1534 ( .A0(n1652), .A1(n1419), .B0(n1648), .B1(n1501), .Y(n1194)
         );
  OAI21XLTS U1535 ( .A0(n1195), .A1(n1194), .B0(n1638), .Y(n1193) );
  OAI31X1TS U1536 ( .A0(n1195), .A1(n1638), .A2(n1194), .B0(n1193), .Y(
        \mult_x_1/n1176 ) );
  OAI22X1TS U1537 ( .A0(n1654), .A1(n1409), .B0(n1518), .B1(n1435), .Y(n1198)
         );
  OAI22X1TS U1538 ( .A0(n1652), .A1(n1413), .B0(n1648), .B1(n1419), .Y(n1197)
         );
  OAI21XLTS U1539 ( .A0(n1198), .A1(n1197), .B0(n1638), .Y(n1196) );
  OAI31X1TS U1540 ( .A0(n1198), .A1(n1638), .A2(n1197), .B0(n1196), .Y(
        \mult_x_1/n1175 ) );
  OAI22X1TS U1541 ( .A0(n1654), .A1(n1427), .B0(n1518), .B1(n1492), .Y(n1201)
         );
  OAI22X1TS U1542 ( .A0(n1652), .A1(n1460), .B0(n1648), .B1(n1461), .Y(n1200)
         );
  OAI21XLTS U1543 ( .A0(n1201), .A1(n1200), .B0(n1638), .Y(n1199) );
  OAI31X1TS U1544 ( .A0(n1201), .A1(n1638), .A2(n1200), .B0(n1199), .Y(
        \mult_x_1/n1165 ) );
  OAI22X1TS U1545 ( .A0(n1654), .A1(n1448), .B0(n1518), .B1(n1449), .Y(n1204)
         );
  OAI22X1TS U1546 ( .A0(n1652), .A1(n1481), .B0(n1648), .B1(n1482), .Y(n1203)
         );
  OAI21XLTS U1547 ( .A0(n1204), .A1(n1203), .B0(n1638), .Y(n1202) );
  OAI31X1TS U1548 ( .A0(n1204), .A1(n1638), .A2(n1203), .B0(n1202), .Y(
        \mult_x_1/n1169 ) );
  OAI22X1TS U1549 ( .A0(n1654), .A1(n1436), .B0(n1518), .B1(n1470), .Y(n1207)
         );
  OAI22X1TS U1550 ( .A0(n1652), .A1(n1468), .B0(n1648), .B1(n1435), .Y(n1206)
         );
  OAI21XLTS U1551 ( .A0(n1207), .A1(n1206), .B0(n1638), .Y(n1205) );
  OAI31X1TS U1552 ( .A0(n1207), .A1(n1638), .A2(n1206), .B0(n1205), .Y(
        \mult_x_1/n1173 ) );
  OAI22X1TS U1553 ( .A0(n1654), .A1(n1414), .B0(n1518), .B1(n1468), .Y(n1210)
         );
  OAI22X1TS U1554 ( .A0(n1652), .A1(n1435), .B0(n1648), .B1(n1413), .Y(n1209)
         );
  OAI21XLTS U1555 ( .A0(n1210), .A1(n1209), .B0(n1638), .Y(n1208) );
  OAI31X1TS U1556 ( .A0(n1210), .A1(n1638), .A2(n1209), .B0(n1208), .Y(
        \mult_x_1/n1174 ) );
  OAI22X1TS U1557 ( .A0(n1654), .A1(n1444), .B0(n1518), .B1(n1482), .Y(n1213)
         );
  OAI22X1TS U1558 ( .A0(n1652), .A1(n1479), .B0(n1648), .B1(n1470), .Y(n1212)
         );
  OAI21XLTS U1559 ( .A0(n1213), .A1(n1212), .B0(n1638), .Y(n1211) );
  OAI31X1TS U1560 ( .A0(n1213), .A1(n1638), .A2(n1212), .B0(n1211), .Y(
        \mult_x_1/n1171 ) );
  OAI22X1TS U1561 ( .A0(n1654), .A1(n1459), .B0(n1518), .B1(n1460), .Y(n1216)
         );
  OAI22X1TS U1562 ( .A0(n1652), .A1(n1461), .B0(n1648), .B1(n1458), .Y(n1215)
         );
  OAI21XLTS U1563 ( .A0(n1216), .A1(n1215), .B0(n1638), .Y(n1214) );
  OAI31X1TS U1564 ( .A0(n1216), .A1(n1638), .A2(n1215), .B0(n1214), .Y(
        \mult_x_1/n1166 ) );
  OAI22X1TS U1565 ( .A0(n1654), .A1(n1469), .B0(n1518), .B1(n1479), .Y(n1219)
         );
  OAI22X1TS U1566 ( .A0(n1652), .A1(n1470), .B0(n1648), .B1(n1468), .Y(n1218)
         );
  OAI21XLTS U1567 ( .A0(n1219), .A1(n1218), .B0(n1638), .Y(n1217) );
  OAI31X1TS U1568 ( .A0(n1219), .A1(n1638), .A2(n1218), .B0(n1217), .Y(
        \mult_x_1/n1172 ) );
  OAI22X1TS U1569 ( .A0(n1654), .A1(n1393), .B0(n1518), .B1(n1461), .Y(n1222)
         );
  OAI22X1TS U1570 ( .A0(n1652), .A1(n1458), .B0(n1648), .B1(n1449), .Y(n1221)
         );
  OAI21XLTS U1571 ( .A0(n1222), .A1(n1221), .B0(n1638), .Y(n1220) );
  OAI31X1TS U1572 ( .A0(n1222), .A1(n1638), .A2(n1221), .B0(n1220), .Y(
        \mult_x_1/n1167 ) );
  OAI22X1TS U1573 ( .A0(n1654), .A1(n1480), .B0(n1518), .B1(n1481), .Y(n1225)
         );
  OAI22X1TS U1574 ( .A0(n1652), .A1(n1482), .B0(n1648), .B1(n1479), .Y(n1224)
         );
  OAI21XLTS U1575 ( .A0(n1225), .A1(n1224), .B0(n1638), .Y(n1223) );
  OAI31X1TS U1576 ( .A0(n1225), .A1(n1638), .A2(n1224), .B0(n1223), .Y(
        \mult_x_1/n1170 ) );
  OAI22X1TS U1577 ( .A0(n1654), .A1(n1418), .B0(n1518), .B1(n1419), .Y(n1228)
         );
  OAI22X1TS U1578 ( .A0(n1652), .A1(n1501), .B0(n1648), .B1(n1506), .Y(n1227)
         );
  OAI21XLTS U1579 ( .A0(n1228), .A1(n1227), .B0(n1638), .Y(n1226) );
  OAI31X1TS U1580 ( .A0(n1228), .A1(n1638), .A2(n1227), .B0(n1226), .Y(
        \mult_x_1/n1177 ) );
  OAI22X1TS U1581 ( .A0(n1654), .A1(n1423), .B0(n1518), .B1(n1458), .Y(n1231)
         );
  OAI22X1TS U1582 ( .A0(n1652), .A1(n1449), .B0(n1648), .B1(n1481), .Y(n1230)
         );
  OAI21XLTS U1583 ( .A0(n1231), .A1(n1230), .B0(n1638), .Y(n1229) );
  OAI31X1TS U1584 ( .A0(n1231), .A1(n1638), .A2(n1230), .B0(n1229), .Y(
        \mult_x_1/n1168 ) );
  OAI22X1TS U1585 ( .A0(n1654), .A1(n1493), .B0(n1518), .B1(n1494), .Y(n1234)
         );
  OAI22X1TS U1586 ( .A0(n1652), .A1(n1495), .B0(n1648), .B1(n1492), .Y(n1233)
         );
  OAI21XLTS U1587 ( .A0(n1234), .A1(n1233), .B0(n1638), .Y(n1232) );
  OAI31X1TS U1588 ( .A0(n1234), .A1(n1638), .A2(n1233), .B0(n1232), .Y(
        \mult_x_1/n1163 ) );
  OAI22X1TS U1589 ( .A0(n1654), .A1(n1401), .B0(n1518), .B1(n1495), .Y(n1237)
         );
  OAI22X1TS U1590 ( .A0(n1652), .A1(n1492), .B0(n1648), .B1(n1460), .Y(n1236)
         );
  OAI21XLTS U1591 ( .A0(n1237), .A1(n1236), .B0(n1638), .Y(n1235) );
  OAI31X1TS U1592 ( .A0(n1237), .A1(n1638), .A2(n1236), .B0(n1235), .Y(
        \mult_x_1/n1164 ) );
  OAI22X1TS U1593 ( .A0(n1654), .A1(n1500), .B0(n1518), .B1(n1501), .Y(n1240)
         );
  OAI22X1TS U1594 ( .A0(n1652), .A1(n1506), .B0(n1648), .B1(n1533), .Y(n1239)
         );
  OAI21XLTS U1595 ( .A0(n1240), .A1(n1239), .B0(n1638), .Y(n1238) );
  OAI31X1TS U1596 ( .A0(n1240), .A1(n1638), .A2(n1239), .B0(n1238), .Y(
        \mult_x_1/n1178 ) );
  OAI22X1TS U1597 ( .A0(n1654), .A1(n1505), .B0(n1518), .B1(n1506), .Y(n1243)
         );
  OAI22X1TS U1598 ( .A0(n1652), .A1(n1533), .B0(n1648), .B1(n1552), .Y(n1242)
         );
  OAI21XLTS U1599 ( .A0(n1243), .A1(n1242), .B0(n1638), .Y(n1241) );
  OAI31X1TS U1600 ( .A0(n1243), .A1(n1638), .A2(n1242), .B0(n1241), .Y(
        \mult_x_1/n1179 ) );
  OAI22X1TS U1601 ( .A0(n1657), .A1(n1561), .B0(n1656), .B1(n1560), .Y(n1246)
         );
  OAI22X1TS U1602 ( .A0(n1322), .A1(n1580), .B0(n1279), .B1(n1650), .Y(n1245)
         );
  OAI21XLTS U1603 ( .A0(n1246), .A1(n1245), .B0(n1674), .Y(n1244) );
  OAI31X1TS U1604 ( .A0(n1246), .A1(n1674), .A2(n1245), .B0(n1244), .Y(
        \mult_x_1/n1191 ) );
  OAI22X1TS U1605 ( .A0(n1657), .A1(n1453), .B0(n1656), .B1(n1475), .Y(n1249)
         );
  OAI22X1TS U1606 ( .A0(n1322), .A1(n1454), .B0(n1279), .B1(n1560), .Y(n1248)
         );
  OAI21XLTS U1607 ( .A0(n1249), .A1(n1248), .B0(n1674), .Y(n1247) );
  OAI31X1TS U1608 ( .A0(n1249), .A1(n1674), .A2(n1248), .B0(n1247), .Y(
        \mult_x_1/n1193 ) );
  OAI22X1TS U1609 ( .A0(n1657), .A1(n1440), .B0(n1656), .B1(n1454), .Y(n1252)
         );
  OAI22X1TS U1610 ( .A0(n1528), .A1(n1560), .B0(n1279), .B1(n1580), .Y(n1251)
         );
  OAI21XLTS U1611 ( .A0(n1252), .A1(n1251), .B0(n1674), .Y(n1250) );
  OAI31X1TS U1612 ( .A0(n1252), .A1(n1674), .A2(n1251), .B0(n1250), .Y(
        \mult_x_1/n1192 ) );
  OAI22X1TS U1613 ( .A0(n1657), .A1(n1397), .B0(n1656), .B1(n1487), .Y(n1255)
         );
  OAI22X1TS U1614 ( .A0(n1322), .A1(n1475), .B0(n1279), .B1(n1454), .Y(n1254)
         );
  OAI21XLTS U1615 ( .A0(n1255), .A1(n1254), .B0(n1674), .Y(n1253) );
  OAI31X1TS U1616 ( .A0(n1255), .A1(n1674), .A2(n1254), .B0(n1253), .Y(
        \mult_x_1/n1194 ) );
  INVX2TS U1617 ( .A(\mult_x_1/n314 ), .Y(n1344) );
  INVX2TS U1618 ( .A(\mult_x_1/n311 ), .Y(n1343) );
  INVX2TS U1619 ( .A(n1259), .Y(Product[56]) );
  OAI22X1TS U1620 ( .A0(n1657), .A1(n1474), .B0(n1656), .B1(n1488), .Y(n1262)
         );
  OAI22X1TS U1621 ( .A0(n1322), .A1(n1487), .B0(n1279), .B1(n1475), .Y(n1261)
         );
  OAI21XLTS U1622 ( .A0(n1262), .A1(n1261), .B0(n1674), .Y(n1260) );
  OAI31X1TS U1623 ( .A0(n1262), .A1(n1674), .A2(n1261), .B0(n1260), .Y(
        \mult_x_1/n1195 ) );
  NOR2XLTS U1624 ( .A(n9), .B(n1263), .Y(\mult_x_1/n759 ) );
  OAI222X1TS U1625 ( .A0(n1646), .A1(n1516), .B0(n1264), .B1(n23), .C0(n1346), 
        .C1(n9), .Y(n1611) );
  AOI21X1TS U1626 ( .A0(A[17]), .A1(\mult_x_1/n759 ), .B0(n1611), .Y(n1632) );
  NAND2X1TS U1627 ( .A(A[17]), .B(n1632), .Y(n1268) );
  OAI22X1TS U1628 ( .A0(n9), .A1(n1645), .B0(n1517), .B1(n1646), .Y(n1266) );
  OAI22X1TS U1629 ( .A0(n29), .A1(n1264), .B0(n23), .B1(n1361), .Y(n1265) );
  NOR2XLTS U1630 ( .A(n1266), .B(n1265), .Y(n1634) );
  INVX2TS U1631 ( .A(n1634), .Y(n1267) );
  OR2X1TS U1632 ( .A(n1268), .B(n1267), .Y(n1631) );
  OAI22X1TS U1633 ( .A0(n1527), .A1(n1646), .B0(n23), .B1(n1645), .Y(n1271) );
  OAI22X1TS U1634 ( .A0(n1554), .A1(n1264), .B0(n29), .B1(n1361), .Y(n1270) );
  OAI21XLTS U1635 ( .A0(n1271), .A1(n1270), .B0(A[17]), .Y(n1269) );
  OAI31X1TS U1636 ( .A0(n1271), .A1(A[17]), .A2(n1270), .B0(n1269), .Y(n1350)
         );
  XNOR2X1TS U1637 ( .A(n1631), .B(n1350), .Y(n1272) );
  XOR2XLTS U1638 ( .A(n1351), .B(n1272), .Y(\mult_x_1/n733 ) );
  OAI22X1TS U1639 ( .A0(n1657), .A1(n1448), .B0(n1656), .B1(n1482), .Y(n1275)
         );
  OAI22X1TS U1640 ( .A0(n1528), .A1(n1481), .B0(n1279), .B1(n1449), .Y(n1274)
         );
  OAI21XLTS U1641 ( .A0(n1275), .A1(n1274), .B0(n1674), .Y(n1273) );
  OAI31X1TS U1642 ( .A0(n1275), .A1(n1674), .A2(n1274), .B0(n1273), .Y(
        \mult_x_1/n1204 ) );
  OAI22X1TS U1643 ( .A0(n1657), .A1(n1393), .B0(n1656), .B1(n1449), .Y(n1278)
         );
  OAI22X1TS U1644 ( .A0(n1322), .A1(n1458), .B0(n1279), .B1(n1461), .Y(n1277)
         );
  OAI21XLTS U1645 ( .A0(n1278), .A1(n1277), .B0(n1674), .Y(n1276) );
  OAI31X1TS U1646 ( .A0(n1278), .A1(n1674), .A2(n1277), .B0(n1276), .Y(
        \mult_x_1/n1202 ) );
  OAI22X1TS U1647 ( .A0(n1657), .A1(n1444), .B0(n1656), .B1(n1470), .Y(n1282)
         );
  OAI22X1TS U1648 ( .A0(n1528), .A1(n1479), .B0(n1279), .B1(n1482), .Y(n1281)
         );
  OAI21XLTS U1649 ( .A0(n1282), .A1(n1281), .B0(n1674), .Y(n1280) );
  OAI31X1TS U1650 ( .A0(n1282), .A1(n1674), .A2(n1281), .B0(n1280), .Y(
        \mult_x_1/n1206 ) );
  OAI22X1TS U1651 ( .A0(n1657), .A1(n1423), .B0(n1656), .B1(n1481), .Y(n1285)
         );
  OAI22X1TS U1652 ( .A0(n1322), .A1(n1449), .B0(n1279), .B1(n1458), .Y(n1284)
         );
  OAI21XLTS U1653 ( .A0(n1285), .A1(n1284), .B0(n1674), .Y(n1283) );
  OAI31X1TS U1654 ( .A0(n1285), .A1(n1674), .A2(n1284), .B0(n1283), .Y(
        \mult_x_1/n1203 ) );
  OAI22X1TS U1655 ( .A0(n1657), .A1(n1469), .B0(n1656), .B1(n1468), .Y(n1288)
         );
  OAI22X1TS U1656 ( .A0(n1528), .A1(n1470), .B0(n1279), .B1(n1479), .Y(n1287)
         );
  OAI21XLTS U1657 ( .A0(n1288), .A1(n1287), .B0(n1674), .Y(n1286) );
  OAI31X1TS U1658 ( .A0(n1288), .A1(n1674), .A2(n1287), .B0(n1286), .Y(
        \mult_x_1/n1207 ) );
  OAI22X1TS U1659 ( .A0(n1657), .A1(n1436), .B0(n1656), .B1(n1435), .Y(n1291)
         );
  OAI22X1TS U1660 ( .A0(n1528), .A1(n1468), .B0(n1279), .B1(n1470), .Y(n1290)
         );
  OAI21XLTS U1661 ( .A0(n1291), .A1(n1290), .B0(n1674), .Y(n1289) );
  OAI31X1TS U1662 ( .A0(n1291), .A1(n1674), .A2(n1290), .B0(n1289), .Y(
        \mult_x_1/n1208 ) );
  OAI22X1TS U1663 ( .A0(n1657), .A1(n1480), .B0(n1656), .B1(n1479), .Y(n1294)
         );
  OAI22X1TS U1664 ( .A0(n1528), .A1(n1482), .B0(n1279), .B1(n1481), .Y(n1293)
         );
  OAI21XLTS U1665 ( .A0(n1294), .A1(n1293), .B0(n1674), .Y(n1292) );
  OAI31X1TS U1666 ( .A0(n1294), .A1(n1674), .A2(n1293), .B0(n1292), .Y(
        \mult_x_1/n1205 ) );
  OAI22X1TS U1667 ( .A0(n1657), .A1(n1431), .B0(n1656), .B1(n1495), .Y(n1297)
         );
  OAI22X1TS U1668 ( .A0(n1322), .A1(n1494), .B0(n1279), .B1(n1488), .Y(n1296)
         );
  OAI21XLTS U1669 ( .A0(n1297), .A1(n1296), .B0(n1674), .Y(n1295) );
  OAI31X1TS U1670 ( .A0(n1297), .A1(n1674), .A2(n1296), .B0(n1295), .Y(
        \mult_x_1/n1197 ) );
  OAI22X1TS U1671 ( .A0(n1657), .A1(n1405), .B0(n1656), .B1(n1501), .Y(n1300)
         );
  OAI22X1TS U1672 ( .A0(n1528), .A1(n1419), .B0(n1279), .B1(n1413), .Y(n1299)
         );
  OAI21XLTS U1673 ( .A0(n1300), .A1(n1299), .B0(n1674), .Y(n1298) );
  OAI31X1TS U1674 ( .A0(n1300), .A1(n1674), .A2(n1299), .B0(n1298), .Y(
        \mult_x_1/n1211 ) );
  OAI22X1TS U1675 ( .A0(n1657), .A1(n1493), .B0(n1656), .B1(n1492), .Y(n1303)
         );
  OAI22X1TS U1676 ( .A0(n1322), .A1(n1495), .B0(n1279), .B1(n1494), .Y(n1302)
         );
  OAI21XLTS U1677 ( .A0(n1303), .A1(n1302), .B0(n1674), .Y(n1301) );
  OAI31X1TS U1678 ( .A0(n1303), .A1(n1674), .A2(n1302), .B0(n1301), .Y(
        \mult_x_1/n1198 ) );
  OAI22X1TS U1679 ( .A0(n1657), .A1(n1409), .B0(n1656), .B1(n1419), .Y(n1306)
         );
  OAI22X1TS U1680 ( .A0(n1528), .A1(n1413), .B0(n1279), .B1(n1435), .Y(n1305)
         );
  OAI21XLTS U1681 ( .A0(n1306), .A1(n1305), .B0(n1674), .Y(n1304) );
  OAI31X1TS U1682 ( .A0(n1306), .A1(n1674), .A2(n1305), .B0(n1304), .Y(
        \mult_x_1/n1210 ) );
  OAI22X1TS U1683 ( .A0(n1657), .A1(n1418), .B0(n1656), .B1(n1506), .Y(n1309)
         );
  OAI22X1TS U1684 ( .A0(n1528), .A1(n1501), .B0(n1279), .B1(n1419), .Y(n1308)
         );
  OAI21XLTS U1685 ( .A0(n1309), .A1(n1308), .B0(n1674), .Y(n1307) );
  OAI31X1TS U1686 ( .A0(n1309), .A1(n1674), .A2(n1308), .B0(n1307), .Y(
        \mult_x_1/n1212 ) );
  OAI22X1TS U1687 ( .A0(n1657), .A1(n1414), .B0(n1656), .B1(n1413), .Y(n1312)
         );
  OAI22X1TS U1688 ( .A0(n1528), .A1(n1435), .B0(n1279), .B1(n1468), .Y(n1311)
         );
  OAI21XLTS U1689 ( .A0(n1312), .A1(n1311), .B0(n1674), .Y(n1310) );
  OAI31X1TS U1690 ( .A0(n1312), .A1(n1674), .A2(n1311), .B0(n1310), .Y(
        \mult_x_1/n1209 ) );
  OAI22X1TS U1691 ( .A0(n1657), .A1(n1427), .B0(n1656), .B1(n1461), .Y(n1315)
         );
  OAI22X1TS U1692 ( .A0(n1322), .A1(n1460), .B0(n1279), .B1(n1492), .Y(n1314)
         );
  OAI21XLTS U1693 ( .A0(n1315), .A1(n1314), .B0(n1674), .Y(n1313) );
  OAI31X1TS U1694 ( .A0(n1315), .A1(n1674), .A2(n1314), .B0(n1313), .Y(
        \mult_x_1/n1200 ) );
  OAI22X1TS U1695 ( .A0(n1657), .A1(n1459), .B0(n1656), .B1(n1458), .Y(n1318)
         );
  OAI22X1TS U1696 ( .A0(n1322), .A1(n1461), .B0(n1279), .B1(n1460), .Y(n1317)
         );
  OAI21XLTS U1697 ( .A0(n1318), .A1(n1317), .B0(n1674), .Y(n1316) );
  OAI31X1TS U1698 ( .A0(n1318), .A1(n1674), .A2(n1317), .B0(n1316), .Y(
        \mult_x_1/n1201 ) );
  OAI22X1TS U1699 ( .A0(n1657), .A1(n1486), .B0(n1656), .B1(n1494), .Y(n1321)
         );
  OAI22X1TS U1700 ( .A0(n1322), .A1(n1488), .B0(n1279), .B1(n1487), .Y(n1320)
         );
  OAI21XLTS U1701 ( .A0(n1321), .A1(n1320), .B0(n1674), .Y(n1319) );
  OAI31X1TS U1702 ( .A0(n1321), .A1(n1674), .A2(n1320), .B0(n1319), .Y(
        \mult_x_1/n1196 ) );
  OAI22X1TS U1703 ( .A0(n1657), .A1(n1401), .B0(n1656), .B1(n1460), .Y(n1325)
         );
  OAI22X1TS U1704 ( .A0(n1322), .A1(n1492), .B0(n1279), .B1(n1495), .Y(n1324)
         );
  OAI21XLTS U1705 ( .A0(n1325), .A1(n1324), .B0(n1674), .Y(n1323) );
  OAI31X1TS U1706 ( .A0(n1325), .A1(n1674), .A2(n1324), .B0(n1323), .Y(
        \mult_x_1/n1199 ) );
  OAI22X1TS U1707 ( .A0(n1657), .A1(n1500), .B0(n1656), .B1(n1533), .Y(n1328)
         );
  OAI22X1TS U1708 ( .A0(n1528), .A1(n1506), .B0(n1279), .B1(n1501), .Y(n1327)
         );
  OAI21XLTS U1709 ( .A0(n1328), .A1(n1327), .B0(n1674), .Y(n1326) );
  OAI31X1TS U1710 ( .A0(n1328), .A1(n1674), .A2(n1327), .B0(n1326), .Y(
        \mult_x_1/n1213 ) );
  OAI22X1TS U1711 ( .A0(n1657), .A1(n1505), .B0(n1656), .B1(n1552), .Y(n1331)
         );
  OAI22X1TS U1712 ( .A0(n1528), .A1(n1533), .B0(n1279), .B1(n1506), .Y(n1330)
         );
  OAI21XLTS U1713 ( .A0(n1331), .A1(n1330), .B0(n1674), .Y(n1329) );
  OAI31X1TS U1714 ( .A0(n1331), .A1(n1674), .A2(n1330), .B0(n1329), .Y(
        \mult_x_1/n1214 ) );
  AOI222XLTS U1715 ( .A0(n1334), .A1(B[31]), .B0(n1333), .B1(n1606), .C0(n1332), .C1(B[30]), .Y(n1335) );
  XOR2XLTS U1716 ( .A(n1674), .B(n1335), .Y(\mult_x_1/n1189 ) );
  OAI22X1TS U1717 ( .A0(n1657), .A1(n1532), .B0(n1656), .B1(n813), .Y(n1338)
         );
  OAI22X1TS U1718 ( .A0(n1528), .A1(n1552), .B0(n1279), .B1(n1533), .Y(n1337)
         );
  OAI21XLTS U1719 ( .A0(n1338), .A1(n1337), .B0(n1674), .Y(n1336) );
  OAI31X1TS U1720 ( .A0(n1338), .A1(n1674), .A2(n1337), .B0(n1336), .Y(
        \mult_x_1/n1215 ) );
  OAI22X1TS U1721 ( .A0(n1654), .A1(n1532), .B0(n1518), .B1(n1533), .Y(n1341)
         );
  OAI22X1TS U1722 ( .A0(n1652), .A1(n1552), .B0(n1648), .B1(n813), .Y(n1340)
         );
  OAI21XLTS U1723 ( .A0(n1341), .A1(n1340), .B0(n1638), .Y(n1339) );
  OAI31X1TS U1724 ( .A0(n1341), .A1(n1638), .A2(n1340), .B0(n1339), .Y(
        \mult_x_1/n1180 ) );
  INVX2TS U1725 ( .A(\mult_x_1/n310 ), .Y(n1375) );
  INVX2TS U1726 ( .A(\mult_x_1/n306 ), .Y(n1374) );
  INVX2TS U1727 ( .A(n1345), .Y(Product[57]) );
  OAI22X1TS U1728 ( .A0(n29), .A1(n1645), .B0(n1646), .B1(n1537), .Y(n1349) );
  OAI22X1TS U1729 ( .A0(n1554), .A1(n1346), .B0(n1264), .B1(n813), .Y(n1348)
         );
  OAI21XLTS U1730 ( .A0(n1349), .A1(n1348), .B0(A[17]), .Y(n1347) );
  OAI31X1TS U1731 ( .A0(n1349), .A1(A[17]), .A2(n1348), .B0(n1347), .Y(n1360)
         );
  AO21XLTS U1732 ( .A0(n1631), .A1(n1351), .B0(n1350), .Y(n1359) );
  OAI31X1TS U1733 ( .A0(n1352), .A1(n1351), .A2(n1672), .B0(n1354), .Y(n1358)
         );
  INVX2TS U1734 ( .A(n1353), .Y(\mult_x_1/n723 ) );
  INVX2TS U1735 ( .A(n1354), .Y(n1357) );
  OAI21XLTS U1736 ( .A0(n1357), .A1(n1672), .B0(n1356), .Y(n1355) );
  OAI31X1TS U1737 ( .A0(n1357), .A1(n1356), .A2(n1672), .B0(n1355), .Y(n1368)
         );
  OAI22X1TS U1738 ( .A0(n1554), .A1(n1645), .B0(n1646), .B1(n1553), .Y(n1364)
         );
  OAI22X1TS U1739 ( .A0(n1361), .A1(n813), .B0(n1264), .B1(n1552), .Y(n1363)
         );
  OAI21XLTS U1740 ( .A0(n1364), .A1(n1363), .B0(A[17]), .Y(n1362) );
  OAI31X1TS U1741 ( .A0(n1364), .A1(A[17]), .A2(n1363), .B0(n1362), .Y(n1366)
         );
  INVX2TS U1742 ( .A(n1365), .Y(\mult_x_1/n712 ) );
  INVX2TS U1743 ( .A(n1369), .Y(\mult_x_1/n713 ) );
  OAI22X1TS U1744 ( .A0(n1554), .A1(n1656), .B0(n1657), .B1(n1553), .Y(n1372)
         );
  OAI22X1TS U1745 ( .A0(n1528), .A1(n813), .B0(n1279), .B1(n1552), .Y(n1371)
         );
  OAI21XLTS U1746 ( .A0(n1372), .A1(n1371), .B0(n1674), .Y(n1370) );
  OAI31X1TS U1747 ( .A0(n1372), .A1(n1674), .A2(n1371), .B0(n1370), .Y(
        \mult_x_1/n1216 ) );
  INVX2TS U1748 ( .A(\mult_x_1/n305 ), .Y(n1391) );
  INVX2TS U1749 ( .A(\mult_x_1/n303 ), .Y(n1390) );
  INVX2TS U1750 ( .A(n1376), .Y(Product[58]) );
  OAI22X1TS U1751 ( .A0(n1660), .A1(n1581), .B0(n1659), .B1(n1580), .Y(n1379)
         );
  OAI22X1TS U1752 ( .A0(n1496), .A1(n1650), .B0(n1507), .B1(n1664), .Y(n1378)
         );
  OAI21XLTS U1753 ( .A0(n1379), .A1(n1378), .B0(n14), .Y(n1377) );
  OAI31X1TS U1754 ( .A0(n1379), .A1(n14), .A2(n1378), .B0(n1377), .Y(
        \mult_x_1/n1225 ) );
  OAI22X1TS U1755 ( .A0(n29), .A1(n1656), .B0(n1657), .B1(n1537), .Y(n1382) );
  OAI22X1TS U1756 ( .A0(n1554), .A1(n1528), .B0(n1279), .B1(n813), .Y(n1381)
         );
  OAI21XLTS U1757 ( .A0(n1382), .A1(n1381), .B0(n1674), .Y(n1380) );
  OAI31X1TS U1758 ( .A0(n1382), .A1(n1674), .A2(n1381), .B0(n1380), .Y(
        \mult_x_1/n1217 ) );
  INVX2TS U1759 ( .A(\mult_x_1/n302 ), .Y(n1571) );
  NOR2XLTS U1760 ( .A(n1580), .B(n1579), .Y(n1384) );
  OAI22X1TS U1761 ( .A0(n1440), .A1(n1592), .B0(n1454), .B1(n1559), .Y(n1383)
         );
  AOI211XLTS U1762 ( .A0(n1584), .A1(B[28]), .B0(n1384), .C0(n1383), .Y(n1568)
         );
  AOI222XLTS U1763 ( .A0(n1387), .A1(n1606), .B0(n1386), .B1(B[31]), .C0(n1385), .C1(B[30]), .Y(n1388) );
  XOR2XLTS U1764 ( .A(n1388), .B(A[29]), .Y(n1567) );
  INVX2TS U1765 ( .A(n1392), .Y(Product[59]) );
  OAI22X1TS U1766 ( .A0(n1660), .A1(n1393), .B0(n1659), .B1(n1449), .Y(n1396)
         );
  OAI22X1TS U1767 ( .A0(n1496), .A1(n1458), .B0(n1507), .B1(n1461), .Y(n1395)
         );
  OAI21XLTS U1768 ( .A0(n1396), .A1(n1395), .B0(n14), .Y(n1394) );
  OAI31X1TS U1769 ( .A0(n1396), .A1(n14), .A2(n1395), .B0(n1394), .Y(
        \mult_x_1/n1237 ) );
  OAI22X1TS U1770 ( .A0(n1660), .A1(n1397), .B0(n1659), .B1(n1487), .Y(n1400)
         );
  OAI22X1TS U1771 ( .A0(n1496), .A1(n1475), .B0(n1507), .B1(n1454), .Y(n1399)
         );
  OAI21XLTS U1772 ( .A0(n1400), .A1(n1399), .B0(n14), .Y(n1398) );
  OAI31X1TS U1773 ( .A0(n1400), .A1(n14), .A2(n1399), .B0(n1398), .Y(
        \mult_x_1/n1229 ) );
  OAI22X1TS U1774 ( .A0(n1660), .A1(n1401), .B0(n1659), .B1(n1460), .Y(n1404)
         );
  OAI22X1TS U1775 ( .A0(n1496), .A1(n1492), .B0(n1507), .B1(n1495), .Y(n1403)
         );
  OAI21XLTS U1776 ( .A0(n1404), .A1(n1403), .B0(n14), .Y(n1402) );
  OAI31X1TS U1777 ( .A0(n1404), .A1(n14), .A2(n1403), .B0(n1402), .Y(
        \mult_x_1/n1234 ) );
  OAI22X1TS U1778 ( .A0(n1660), .A1(n1405), .B0(n1659), .B1(n1501), .Y(n1408)
         );
  OAI22X1TS U1779 ( .A0(n1496), .A1(n1419), .B0(n1507), .B1(n1413), .Y(n1407)
         );
  OAI21XLTS U1780 ( .A0(n1408), .A1(n1407), .B0(n14), .Y(n1406) );
  OAI31X1TS U1781 ( .A0(n1408), .A1(n14), .A2(n1407), .B0(n1406), .Y(
        \mult_x_1/n1246 ) );
  OAI22X1TS U1782 ( .A0(n1660), .A1(n1409), .B0(n1659), .B1(n1419), .Y(n1412)
         );
  OAI22X1TS U1783 ( .A0(n1496), .A1(n1413), .B0(n1507), .B1(n1435), .Y(n1411)
         );
  OAI21XLTS U1784 ( .A0(n1412), .A1(n1411), .B0(n14), .Y(n1410) );
  OAI31X1TS U1785 ( .A0(n1412), .A1(n14), .A2(n1411), .B0(n1410), .Y(
        \mult_x_1/n1245 ) );
  OAI22X1TS U1786 ( .A0(n1660), .A1(n1414), .B0(n1659), .B1(n1413), .Y(n1417)
         );
  OAI22X1TS U1787 ( .A0(n1496), .A1(n1435), .B0(n1507), .B1(n1468), .Y(n1416)
         );
  OAI21XLTS U1788 ( .A0(n1417), .A1(n1416), .B0(n14), .Y(n1415) );
  OAI31X1TS U1789 ( .A0(n1417), .A1(n14), .A2(n1416), .B0(n1415), .Y(
        \mult_x_1/n1244 ) );
  OAI22X1TS U1790 ( .A0(n1660), .A1(n1418), .B0(n1659), .B1(n1506), .Y(n1422)
         );
  OAI22X1TS U1791 ( .A0(n1496), .A1(n1501), .B0(n1507), .B1(n1419), .Y(n1421)
         );
  OAI21XLTS U1792 ( .A0(n1422), .A1(n1421), .B0(n14), .Y(n1420) );
  OAI31X1TS U1793 ( .A0(n1422), .A1(n14), .A2(n1421), .B0(n1420), .Y(
        \mult_x_1/n1247 ) );
  OAI22X1TS U1794 ( .A0(n1660), .A1(n1423), .B0(n1659), .B1(n1481), .Y(n1426)
         );
  OAI22X1TS U1795 ( .A0(n1496), .A1(n1449), .B0(n1507), .B1(n1458), .Y(n1425)
         );
  OAI21XLTS U1796 ( .A0(n1426), .A1(n1425), .B0(n14), .Y(n1424) );
  OAI31X1TS U1797 ( .A0(n1426), .A1(n14), .A2(n1425), .B0(n1424), .Y(
        \mult_x_1/n1238 ) );
  OAI22X1TS U1798 ( .A0(n1660), .A1(n1427), .B0(n1659), .B1(n1461), .Y(n1430)
         );
  OAI22X1TS U1799 ( .A0(n1496), .A1(n1460), .B0(n1507), .B1(n1492), .Y(n1429)
         );
  OAI21XLTS U1800 ( .A0(n1430), .A1(n1429), .B0(n14), .Y(n1428) );
  OAI31X1TS U1801 ( .A0(n1430), .A1(n14), .A2(n1429), .B0(n1428), .Y(
        \mult_x_1/n1235 ) );
  OAI22X1TS U1802 ( .A0(n1660), .A1(n1431), .B0(n1659), .B1(n1495), .Y(n1434)
         );
  OAI22X1TS U1803 ( .A0(n1496), .A1(n1494), .B0(n1507), .B1(n1488), .Y(n1433)
         );
  OAI21XLTS U1804 ( .A0(n1434), .A1(n1433), .B0(n14), .Y(n1432) );
  OAI31X1TS U1805 ( .A0(n1434), .A1(n14), .A2(n1433), .B0(n1432), .Y(
        \mult_x_1/n1232 ) );
  OAI22X1TS U1806 ( .A0(n1660), .A1(n1436), .B0(n1659), .B1(n1435), .Y(n1439)
         );
  OAI22X1TS U1807 ( .A0(n1496), .A1(n1468), .B0(n1507), .B1(n1470), .Y(n1438)
         );
  OAI21XLTS U1808 ( .A0(n1439), .A1(n1438), .B0(n14), .Y(n1437) );
  OAI31X1TS U1809 ( .A0(n1439), .A1(n14), .A2(n1438), .B0(n1437), .Y(
        \mult_x_1/n1243 ) );
  OAI22X1TS U1810 ( .A0(n1660), .A1(n1440), .B0(n1659), .B1(n1454), .Y(n1443)
         );
  OAI22X1TS U1811 ( .A0(n1496), .A1(n1560), .B0(n1507), .B1(n1580), .Y(n1442)
         );
  OAI21XLTS U1812 ( .A0(n1443), .A1(n1442), .B0(n14), .Y(n1441) );
  OAI31X1TS U1813 ( .A0(n1443), .A1(n14), .A2(n1442), .B0(n1441), .Y(
        \mult_x_1/n1227 ) );
  OAI22X1TS U1814 ( .A0(n1660), .A1(n1444), .B0(n1659), .B1(n1470), .Y(n1447)
         );
  OAI22X1TS U1815 ( .A0(n1496), .A1(n1479), .B0(n1507), .B1(n1482), .Y(n1446)
         );
  OAI21XLTS U1816 ( .A0(n1447), .A1(n1446), .B0(n14), .Y(n1445) );
  OAI31X1TS U1817 ( .A0(n1447), .A1(n14), .A2(n1446), .B0(n1445), .Y(
        \mult_x_1/n1241 ) );
  OAI22X1TS U1818 ( .A0(n1660), .A1(n1448), .B0(n1659), .B1(n1482), .Y(n1452)
         );
  OAI22X1TS U1819 ( .A0(n1496), .A1(n1481), .B0(n1507), .B1(n1449), .Y(n1451)
         );
  OAI21XLTS U1820 ( .A0(n1452), .A1(n1451), .B0(n14), .Y(n1450) );
  OAI31X1TS U1821 ( .A0(n1452), .A1(n14), .A2(n1451), .B0(n1450), .Y(
        \mult_x_1/n1239 ) );
  OAI22X1TS U1822 ( .A0(n1660), .A1(n1453), .B0(n1659), .B1(n1475), .Y(n1457)
         );
  OAI22X1TS U1823 ( .A0(n1496), .A1(n1454), .B0(n1507), .B1(n1560), .Y(n1456)
         );
  OAI21XLTS U1824 ( .A0(n1457), .A1(n1456), .B0(n14), .Y(n1455) );
  OAI31X1TS U1825 ( .A0(n1457), .A1(n14), .A2(n1456), .B0(n1455), .Y(
        \mult_x_1/n1228 ) );
  OAI22X1TS U1826 ( .A0(n1660), .A1(n1459), .B0(n1659), .B1(n1458), .Y(n1464)
         );
  OAI22X1TS U1827 ( .A0(n1496), .A1(n1461), .B0(n1507), .B1(n1460), .Y(n1463)
         );
  OAI21XLTS U1828 ( .A0(n1464), .A1(n1463), .B0(n14), .Y(n1462) );
  OAI31X1TS U1829 ( .A0(n1464), .A1(n14), .A2(n1463), .B0(n1462), .Y(
        \mult_x_1/n1236 ) );
  OAI22X1TS U1830 ( .A0(n1660), .A1(n1561), .B0(n1659), .B1(n1560), .Y(n1467)
         );
  OAI22X1TS U1831 ( .A0(n1496), .A1(n1580), .B0(n1507), .B1(n1650), .Y(n1466)
         );
  OAI21XLTS U1832 ( .A0(n1467), .A1(n1466), .B0(n14), .Y(n1465) );
  OAI31X1TS U1833 ( .A0(n1467), .A1(n14), .A2(n1466), .B0(n1465), .Y(
        \mult_x_1/n1226 ) );
  OAI22X1TS U1834 ( .A0(n1660), .A1(n1469), .B0(n1659), .B1(n1468), .Y(n1473)
         );
  OAI22X1TS U1835 ( .A0(n1496), .A1(n1470), .B0(n1507), .B1(n1479), .Y(n1472)
         );
  OAI21XLTS U1836 ( .A0(n1473), .A1(n1472), .B0(n14), .Y(n1471) );
  OAI31X1TS U1837 ( .A0(n1473), .A1(n14), .A2(n1472), .B0(n1471), .Y(
        \mult_x_1/n1242 ) );
  OAI22X1TS U1838 ( .A0(n1660), .A1(n1474), .B0(n1659), .B1(n1488), .Y(n1478)
         );
  OAI22X1TS U1839 ( .A0(n1496), .A1(n1487), .B0(n1507), .B1(n1475), .Y(n1477)
         );
  OAI21XLTS U1840 ( .A0(n1478), .A1(n1477), .B0(n14), .Y(n1476) );
  OAI31X1TS U1841 ( .A0(n1478), .A1(n14), .A2(n1477), .B0(n1476), .Y(
        \mult_x_1/n1230 ) );
  OAI22X1TS U1842 ( .A0(n1660), .A1(n1480), .B0(n1659), .B1(n1479), .Y(n1485)
         );
  OAI22X1TS U1843 ( .A0(n1496), .A1(n1482), .B0(n1507), .B1(n1481), .Y(n1484)
         );
  OAI21XLTS U1844 ( .A0(n1485), .A1(n1484), .B0(n14), .Y(n1483) );
  OAI31X1TS U1845 ( .A0(n1485), .A1(n14), .A2(n1484), .B0(n1483), .Y(
        \mult_x_1/n1240 ) );
  OAI22X1TS U1846 ( .A0(n1660), .A1(n1486), .B0(n1659), .B1(n1494), .Y(n1491)
         );
  OAI22X1TS U1847 ( .A0(n1496), .A1(n1488), .B0(n1507), .B1(n1487), .Y(n1490)
         );
  OAI21XLTS U1848 ( .A0(n1491), .A1(n1490), .B0(n14), .Y(n1489) );
  OAI31X1TS U1849 ( .A0(n1491), .A1(n14), .A2(n1490), .B0(n1489), .Y(
        \mult_x_1/n1231 ) );
  OAI22X1TS U1850 ( .A0(n1660), .A1(n1493), .B0(n1659), .B1(n1492), .Y(n1499)
         );
  OAI22X1TS U1851 ( .A0(n1496), .A1(n1495), .B0(n1507), .B1(n1494), .Y(n1498)
         );
  OAI21XLTS U1852 ( .A0(n1499), .A1(n1498), .B0(n14), .Y(n1497) );
  OAI31X1TS U1853 ( .A0(n1499), .A1(n14), .A2(n1498), .B0(n1497), .Y(
        \mult_x_1/n1233 ) );
  OAI22X1TS U1854 ( .A0(n1660), .A1(n1500), .B0(n1659), .B1(n1533), .Y(n1504)
         );
  OAI22X1TS U1855 ( .A0(n1496), .A1(n1506), .B0(n1507), .B1(n1501), .Y(n1503)
         );
  OAI21XLTS U1856 ( .A0(n1504), .A1(n1503), .B0(n14), .Y(n1502) );
  OAI31X1TS U1857 ( .A0(n1504), .A1(n14), .A2(n1503), .B0(n1502), .Y(
        \mult_x_1/n1248 ) );
  OAI22X1TS U1858 ( .A0(n1660), .A1(n1505), .B0(n1659), .B1(n1552), .Y(n1510)
         );
  OAI22X1TS U1859 ( .A0(n1496), .A1(n1533), .B0(n1507), .B1(n1506), .Y(n1509)
         );
  OAI21XLTS U1860 ( .A0(n1510), .A1(n1509), .B0(n14), .Y(n1508) );
  OAI31X1TS U1861 ( .A0(n1510), .A1(n14), .A2(n1509), .B0(n1508), .Y(
        \mult_x_1/n1249 ) );
  AOI222XLTS U1862 ( .A0(n1513), .A1(n1606), .B0(n1512), .B1(B[31]), .C0(n1511), .C1(B[30]), .Y(n1514) );
  XOR2XLTS U1863 ( .A(n14), .B(n1514), .Y(\mult_x_1/n1224 ) );
  NOR2XLTS U1864 ( .A(n9), .B(n1515), .Y(\mult_x_1/n795 ) );
  OAI222X1TS U1865 ( .A0(n1654), .A1(n1516), .B0(n1518), .B1(n23), .C0(n1652), 
        .C1(n9), .Y(n1612) );
  AOI21X1TS U1866 ( .A0(A[11]), .A1(\mult_x_1/n795 ), .B0(n1612), .Y(n1636) );
  INVX2TS U1867 ( .A(n1636), .Y(n1522) );
  OAI22X1TS U1868 ( .A0(n29), .A1(n1518), .B0(n1517), .B1(n1654), .Y(n1520) );
  OAI22X1TS U1869 ( .A0(n23), .A1(n1652), .B0(n9), .B1(n1648), .Y(n1519) );
  NOR2XLTS U1870 ( .A(n1520), .B(n1519), .Y(n1639) );
  NAND2X1TS U1871 ( .A(A[11]), .B(n1639), .Y(n1521) );
  OR2X1TS U1872 ( .A(n1522), .B(n1521), .Y(n1635) );
  OAI22X1TS U1873 ( .A0(n1554), .A1(n1518), .B0(n1527), .B1(n1654), .Y(n1525)
         );
  OAI22X1TS U1874 ( .A0(n29), .A1(n1652), .B0(n23), .B1(n1648), .Y(n1524) );
  OAI21XLTS U1875 ( .A0(n1525), .A1(n1524), .B0(A[11]), .Y(n1523) );
  OAI31X1TS U1876 ( .A0(n1525), .A1(A[11]), .A2(n1524), .B0(n1523), .Y(n1541)
         );
  XNOR2X1TS U1877 ( .A(n1635), .B(n1541), .Y(n1526) );
  XOR2XLTS U1878 ( .A(n1542), .B(n1526), .Y(\mult_x_1/n778 ) );
  OAI22X1TS U1879 ( .A0(n1527), .A1(n1657), .B0(n23), .B1(n1656), .Y(n1531) );
  OAI22X1TS U1880 ( .A0(n1554), .A1(n1279), .B0(n29), .B1(n1528), .Y(n1530) );
  OAI21XLTS U1881 ( .A0(n1531), .A1(n1530), .B0(n1674), .Y(n1529) );
  OAI31X1TS U1882 ( .A0(n1531), .A1(n1674), .A2(n1530), .B0(n1529), .Y(
        \mult_x_1/n1218 ) );
  OAI22X1TS U1883 ( .A0(n1660), .A1(n1532), .B0(n1659), .B1(n813), .Y(n1536)
         );
  OAI22X1TS U1884 ( .A0(n1496), .A1(n1552), .B0(n1507), .B1(n1533), .Y(n1535)
         );
  OAI21XLTS U1885 ( .A0(n1536), .A1(n1535), .B0(n14), .Y(n1534) );
  OAI31X1TS U1886 ( .A0(n1536), .A1(n14), .A2(n1535), .B0(n1534), .Y(
        \mult_x_1/n1250 ) );
  OAI22X1TS U1887 ( .A0(n1654), .A1(n1537), .B0(n1518), .B1(n813), .Y(n1540)
         );
  OAI22X1TS U1888 ( .A0(n1554), .A1(n1652), .B0(n29), .B1(n1648), .Y(n1539) );
  OAI21XLTS U1889 ( .A0(n1540), .A1(n1539), .B0(A[11]), .Y(n1538) );
  OAI31X1TS U1890 ( .A0(n1540), .A1(A[11]), .A2(n1539), .B0(n1538), .Y(n1551)
         );
  AO21XLTS U1891 ( .A0(n1635), .A1(n1542), .B0(n1541), .Y(n1550) );
  OAI31X1TS U1892 ( .A0(n1543), .A1(n1542), .A2(n1673), .B0(n1545), .Y(n1549)
         );
  INVX2TS U1893 ( .A(n1544), .Y(\mult_x_1/n771 ) );
  INVX2TS U1894 ( .A(n1545), .Y(n1548) );
  OAI21XLTS U1895 ( .A0(n1548), .A1(n1673), .B0(n1547), .Y(n1546) );
  OAI31X1TS U1896 ( .A0(n1548), .A1(n1547), .A2(n1673), .B0(n1546), .Y(n1575)
         );
  OAI22X1TS U1897 ( .A0(n1654), .A1(n1553), .B0(n1518), .B1(n1552), .Y(n1557)
         );
  OAI22X1TS U1898 ( .A0(n1554), .A1(n1648), .B0(n1652), .B1(n813), .Y(n1556)
         );
  OAI21XLTS U1899 ( .A0(n1557), .A1(n1556), .B0(A[11]), .Y(n1555) );
  OAI31X1TS U1900 ( .A0(n1557), .A1(A[11]), .A2(n1556), .B0(n1555), .Y(n1573)
         );
  INVX2TS U1901 ( .A(n1558), .Y(\mult_x_1/n763 ) );
  NOR2XLTS U1902 ( .A(n1650), .B(n1579), .Y(n1563) );
  OAI22X1TS U1903 ( .A0(n1561), .A1(n1663), .B0(n1560), .B1(n1559), .Y(n1562)
         );
  AOI211XLTS U1904 ( .A0(n1584), .A1(B[29]), .B0(n1563), .C0(n1562), .Y(n1578)
         );
  OAI22X1TS U1905 ( .A0(n1565), .A1(n1662), .B0(n1564), .B1(n1664), .Y(n1566)
         );
  XOR2XLTS U1906 ( .A(n1625), .B(n1566), .Y(n1577) );
  INVX2TS U1907 ( .A(n1572), .Y(Product[60]) );
  INVX2TS U1908 ( .A(n1576), .Y(\mult_x_1/n764 ) );
  INVX2TS U1909 ( .A(\mult_x_1/n297 ), .Y(n1590) );
  NOR2XLTS U1910 ( .A(n1664), .B(n1579), .Y(n1583) );
  OAI22X1TS U1911 ( .A0(n1581), .A1(n1663), .B0(n1580), .B1(n1559), .Y(n1582)
         );
  AOI211XLTS U1912 ( .A0(n1584), .A1(B[30]), .B0(n1583), .C0(n1582), .Y(n1589)
         );
  INVX2TS U1913 ( .A(n1588), .Y(Product[61]) );
  OAI222X1TS U1914 ( .A0(n1653), .A1(n1592), .B0(n1591), .B1(n1664), .C0(n1650), .C1(n1559), .Y(n1667) );
  INVX2TS U1915 ( .A(n1596), .Y(Product[62]) );
  INVX2TS U1916 ( .A(n1600), .Y(\mult_x_1/n796 ) );
  OAI22X1TS U1917 ( .A0(n1602), .A1(n1662), .B0(n1601), .B1(n1664), .Y(n1603)
         );
  XOR2XLTS U1918 ( .A(A[26]), .B(n1603), .Y(\mult_x_1/n978 ) );
  AOI222XLTS U1919 ( .A0(n1607), .A1(n1606), .B0(n1605), .B1(B[31]), .C0(n1604), .C1(B[30]), .Y(n1608) );
  XOR2XLTS U1920 ( .A(n539), .B(n1608), .Y(\mult_x_1/n1084 ) );
  AOI31XLTS U1921 ( .A0(A[23]), .A1(\mult_x_1/n705 ), .A2(n1610), .B0(n1609), 
        .Y(\mult_x_1/n694 ) );
  AOI31XLTS U1922 ( .A0(A[17]), .A1(\mult_x_1/n759 ), .A2(n1611), .B0(n1632), 
        .Y(\mult_x_1/n751 ) );
  AOI31XLTS U1923 ( .A0(A[11]), .A1(\mult_x_1/n795 ), .A2(n1612), .B0(n1636), 
        .Y(\mult_x_1/n790 ) );
  OA21XLTS U1924 ( .A0(n1615), .A1(n1614), .B0(n1613), .Y(Product[3]) );
  NAND2X1TS U1925 ( .A(n1616), .B(Product[0]), .Y(n1618) );
  OA21XLTS U1926 ( .A0(n1619), .A1(n1618), .B0(n1617), .Y(Product[1]) );
  OAI31X1TS U1927 ( .A0(n1623), .A1(n1626), .A2(n1625), .B0(n1622), .Y(n1624)
         );
  AOI21X1TS U1928 ( .A0(n1626), .A1(n1625), .B0(n1624), .Y(\mult_x_1/n605 ) );
  XOR2XLTS U1929 ( .A(n1628), .B(n1627), .Y(n1629) );
  XOR2XLTS U1930 ( .A(n1630), .B(n1629), .Y(\mult_x_1/n670 ) );
  OAI31X1TS U1931 ( .A0(n1632), .A1(n1634), .A2(n539), .B0(n1631), .Y(n1633)
         );
  AOI21X1TS U1932 ( .A0(n1634), .A1(n539), .B0(n1633), .Y(\mult_x_1/n743 ) );
  OAI31X1TS U1933 ( .A0(n1636), .A1(n1639), .A2(n1638), .B0(n1635), .Y(n1637)
         );
  AOI21X1TS U1934 ( .A0(n1639), .A1(n1638), .B0(n1637), .Y(\mult_x_1/n785 ) );
  OAI22X1TS U1935 ( .A0(n723), .A1(n1662), .B0(n1640), .B1(n1664), .Y(n1641)
         );
  XOR2XLTS U1936 ( .A(A[23]), .B(n1641), .Y(\mult_x_1/n1013 ) );
  OAI222X1TS U1937 ( .A0(n723), .A1(n1653), .B0(n1643), .B1(n1664), .C0(n1642), 
        .C1(n1650), .Y(n1644) );
  XOR2XLTS U1938 ( .A(A[23]), .B(n1644), .Y(\mult_x_1/n1014 ) );
  OAI22X1TS U1939 ( .A0(n1646), .A1(n1662), .B0(n1645), .B1(n1664), .Y(n1647)
         );
  XOR2XLTS U1940 ( .A(A[17]), .B(n1647), .Y(\mult_x_1/n1083 ) );
  OAI22X1TS U1941 ( .A0(n1654), .A1(n1662), .B0(n1648), .B1(n1664), .Y(n1649)
         );
  XOR2XLTS U1942 ( .A(A[11]), .B(n1649), .Y(\mult_x_1/n1153 ) );
  OAI222X1TS U1943 ( .A0(n1654), .A1(n1653), .B0(n1652), .B1(n1664), .C0(n1651), .C1(n1650), .Y(n1655) );
  XOR2XLTS U1944 ( .A(A[11]), .B(n1655), .Y(\mult_x_1/n1154 ) );
  OAI22X1TS U1945 ( .A0(n1657), .A1(n1662), .B0(n1656), .B1(n1664), .Y(n1658)
         );
  XOR2XLTS U1946 ( .A(A[8]), .B(n1658), .Y(\mult_x_1/n1188 ) );
  OAI22X1TS U1947 ( .A0(n1660), .A1(n1662), .B0(n1659), .B1(n1664), .Y(n1661)
         );
  XOR2XLTS U1948 ( .A(A[5]), .B(n1661), .Y(\mult_x_1/n1223 ) );
  OAI22X1TS U1949 ( .A0(n1664), .A1(n1559), .B0(n1663), .B1(n1662), .Y(n1670)
         );
  XOR2XLTS U1950 ( .A(n1668), .B(n1667), .Y(n1669) );
  XOR2XLTS U1951 ( .A(n1670), .B(n1669), .Y(Product[63]) );
endmodule


module RF ( clk, data_in, data_outA, data_outB, WA, RAA, RAB, enable );
  input [31:0] data_in;
  output [31:0] data_outA;
  output [31:0] data_outB;
  input [5:0] WA;
  input [5:0] RAA;
  input [5:0] RAB;
  input [2:0] enable;
  input clk;
  wire   \Mem[35][31] , \Mem[35][30] , \Mem[35][29] , \Mem[35][28] ,
         \Mem[35][27] , \Mem[35][26] , \Mem[35][25] , \Mem[35][24] ,
         \Mem[35][23] , \Mem[35][22] , \Mem[35][21] , \Mem[35][20] ,
         \Mem[35][19] , \Mem[35][18] , \Mem[35][17] , \Mem[35][16] ,
         \Mem[35][15] , \Mem[35][14] , \Mem[35][13] , \Mem[35][12] ,
         \Mem[35][11] , \Mem[35][10] , \Mem[35][9] , \Mem[35][8] ,
         \Mem[35][7] , \Mem[35][6] , \Mem[35][5] , \Mem[35][4] , \Mem[35][3] ,
         \Mem[35][2] , \Mem[35][1] , \Mem[35][0] , \Mem[34][31] ,
         \Mem[34][30] , \Mem[34][29] , \Mem[34][28] , \Mem[34][27] ,
         \Mem[34][26] , \Mem[34][25] , \Mem[34][24] , \Mem[34][23] ,
         \Mem[34][22] , \Mem[34][21] , \Mem[34][20] , \Mem[34][19] ,
         \Mem[34][18] , \Mem[34][17] , \Mem[34][16] , \Mem[34][15] ,
         \Mem[34][14] , \Mem[34][13] , \Mem[34][12] , \Mem[34][11] ,
         \Mem[34][10] , \Mem[34][9] , \Mem[34][8] , \Mem[34][7] , \Mem[34][6] ,
         \Mem[34][5] , \Mem[34][4] , \Mem[34][3] , \Mem[34][2] , \Mem[34][1] ,
         \Mem[34][0] , \Mem[33][31] , \Mem[33][30] , \Mem[33][29] ,
         \Mem[33][28] , \Mem[33][27] , \Mem[33][26] , \Mem[33][25] ,
         \Mem[33][24] , \Mem[33][23] , \Mem[33][22] , \Mem[33][21] ,
         \Mem[33][20] , \Mem[33][19] , \Mem[33][18] , \Mem[33][17] ,
         \Mem[33][16] , \Mem[33][15] , \Mem[33][14] , \Mem[33][13] ,
         \Mem[33][12] , \Mem[33][11] , \Mem[33][10] , \Mem[33][9] ,
         \Mem[33][8] , \Mem[33][7] , \Mem[33][6] , \Mem[33][5] , \Mem[33][4] ,
         \Mem[33][3] , \Mem[33][2] , \Mem[33][1] , \Mem[33][0] , \Mem[32][31] ,
         \Mem[32][30] , \Mem[32][29] , \Mem[32][28] , \Mem[32][27] ,
         \Mem[32][26] , \Mem[32][25] , \Mem[32][24] , \Mem[32][23] ,
         \Mem[32][22] , \Mem[32][21] , \Mem[32][20] , \Mem[32][19] ,
         \Mem[32][18] , \Mem[32][17] , \Mem[32][16] , \Mem[32][15] ,
         \Mem[32][14] , \Mem[32][13] , \Mem[32][12] , \Mem[32][11] ,
         \Mem[32][10] , \Mem[32][9] , \Mem[32][8] , \Mem[32][7] , \Mem[32][6] ,
         \Mem[32][5] , \Mem[32][4] , \Mem[32][3] , \Mem[32][2] , \Mem[32][1] ,
         \Mem[32][0] , N63, N64, N65, N66, N67, N68, N69, N71, N73, N75, N77,
         N79, N81, N83, N85, N87, N89, N91, N92, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N162, N1928, N1929, N1930, N1931, N1932, N1933, N1934,
         N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944,
         N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953, N1954,
         N1955, N1956, N1957, N1958, N1959, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526;
  assign N162 = enable[0];

  TLATXLTS \data_outB_reg[22]  ( .G(n526), .D(N102), .Q(data_outB[22]) );
  TLATXLTS \data_outB_reg[20]  ( .G(n526), .D(N104), .Q(data_outB[20]) );
  TLATXLTS \data_outB_reg[18]  ( .G(n526), .D(N106), .Q(data_outB[18]) );
  TLATXLTS \data_outB_reg[16]  ( .G(n526), .D(N108), .Q(data_outB[16]) );
  TLATXLTS \data_outB_reg[14]  ( .G(n526), .D(N110), .Q(data_outB[14]) );
  TLATXLTS \data_outB_reg[12]  ( .G(n526), .D(N112), .Q(data_outB[12]) );
  TLATXLTS \data_outB_reg[10]  ( .G(n526), .D(N114), .Q(data_outB[10]) );
  TLATXLTS \data_outB_reg[8]  ( .G(n526), .D(N116), .Q(data_outB[8]) );
  TLATXLTS \data_outB_reg[31]  ( .G(n526), .D(n512), .Q(data_outB[31]) );
  TLATXLTS \data_outB_reg[30]  ( .G(n526), .D(n511), .Q(data_outB[30]) );
  TLATXLTS \data_outB_reg[29]  ( .G(n526), .D(N95), .Q(data_outB[29]) );
  TLATXLTS \data_outB_reg[28]  ( .G(n526), .D(N96), .Q(data_outB[28]) );
  TLATXLTS \data_outB_reg[27]  ( .G(n526), .D(N97), .Q(data_outB[27]) );
  TLATXLTS \data_outB_reg[26]  ( .G(n526), .D(N98), .Q(data_outB[26]) );
  TLATXLTS \data_outB_reg[25]  ( .G(n526), .D(N99), .Q(data_outB[25]) );
  TLATXLTS \data_outB_reg[24]  ( .G(n526), .D(N100), .Q(data_outB[24]) );
  TLATXLTS \data_outB_reg[23]  ( .G(n526), .D(N101), .Q(data_outB[23]) );
  TLATXLTS \data_outB_reg[21]  ( .G(n526), .D(N103), .Q(data_outB[21]) );
  TLATXLTS \data_outB_reg[19]  ( .G(n526), .D(N105), .Q(data_outB[19]) );
  TLATXLTS \data_outB_reg[17]  ( .G(n526), .D(N107), .Q(data_outB[17]) );
  TLATXLTS \data_outB_reg[15]  ( .G(n526), .D(N109), .Q(data_outB[15]) );
  TLATXLTS \data_outB_reg[13]  ( .G(n526), .D(N111), .Q(data_outB[13]) );
  TLATXLTS \data_outB_reg[11]  ( .G(n526), .D(N113), .Q(data_outB[11]) );
  TLATXLTS \data_outB_reg[9]  ( .G(n526), .D(N115), .Q(data_outB[9]) );
  TLATXLTS \data_outB_reg[7]  ( .G(n526), .D(N117), .Q(data_outB[7]) );
  TLATXLTS \data_outB_reg[6]  ( .G(n526), .D(N118), .Q(data_outB[6]) );
  TLATXLTS \data_outB_reg[5]  ( .G(n526), .D(N119), .Q(data_outB[5]) );
  TLATXLTS \data_outB_reg[4]  ( .G(n526), .D(N120), .Q(data_outB[4]) );
  TLATXLTS \data_outB_reg[3]  ( .G(n526), .D(N121), .Q(data_outB[3]) );
  TLATXLTS \data_outB_reg[2]  ( .G(n526), .D(N122), .Q(data_outB[2]) );
  TLATXLTS \data_outB_reg[1]  ( .G(n526), .D(N123), .Q(data_outB[1]) );
  TLATXLTS \data_outB_reg[0]  ( .G(n526), .D(N124), .Q(data_outB[0]) );
  DFFQX1TS \Mem_reg[35][31]  ( .D(N1959), .CK(clk), .Q(\Mem[35][31] ) );
  DFFQX1TS \Mem_reg[35][30]  ( .D(N1958), .CK(clk), .Q(\Mem[35][30] ) );
  DFFQX1TS \Mem_reg[35][29]  ( .D(N1957), .CK(clk), .Q(\Mem[35][29] ) );
  DFFQX1TS \Mem_reg[35][28]  ( .D(N1956), .CK(clk), .Q(\Mem[35][28] ) );
  DFFQX1TS \Mem_reg[35][27]  ( .D(N1955), .CK(clk), .Q(\Mem[35][27] ) );
  DFFQX1TS \Mem_reg[35][26]  ( .D(N1954), .CK(clk), .Q(\Mem[35][26] ) );
  DFFQX1TS \Mem_reg[35][25]  ( .D(N1953), .CK(clk), .Q(\Mem[35][25] ) );
  DFFQX1TS \Mem_reg[35][24]  ( .D(N1952), .CK(clk), .Q(\Mem[35][24] ) );
  DFFQX1TS \Mem_reg[35][23]  ( .D(N1951), .CK(clk), .Q(\Mem[35][23] ) );
  DFFQX1TS \Mem_reg[35][22]  ( .D(N1950), .CK(clk), .Q(\Mem[35][22] ) );
  DFFQX1TS \Mem_reg[35][21]  ( .D(N1949), .CK(clk), .Q(\Mem[35][21] ) );
  DFFQX1TS \Mem_reg[35][20]  ( .D(N1948), .CK(clk), .Q(\Mem[35][20] ) );
  DFFQX1TS \Mem_reg[35][19]  ( .D(N1947), .CK(clk), .Q(\Mem[35][19] ) );
  DFFQX1TS \Mem_reg[35][18]  ( .D(N1946), .CK(clk), .Q(\Mem[35][18] ) );
  DFFQX1TS \Mem_reg[35][17]  ( .D(N1945), .CK(clk), .Q(\Mem[35][17] ) );
  DFFQX1TS \Mem_reg[35][16]  ( .D(N1944), .CK(clk), .Q(\Mem[35][16] ) );
  DFFQX1TS \Mem_reg[35][15]  ( .D(N1943), .CK(clk), .Q(\Mem[35][15] ) );
  DFFQX1TS \Mem_reg[35][14]  ( .D(N1942), .CK(clk), .Q(\Mem[35][14] ) );
  DFFQX1TS \Mem_reg[35][13]  ( .D(N1941), .CK(clk), .Q(\Mem[35][13] ) );
  DFFQX1TS \Mem_reg[35][12]  ( .D(N1940), .CK(clk), .Q(\Mem[35][12] ) );
  DFFQX1TS \Mem_reg[35][11]  ( .D(N1939), .CK(clk), .Q(\Mem[35][11] ) );
  DFFQX1TS \Mem_reg[35][10]  ( .D(N1938), .CK(clk), .Q(\Mem[35][10] ) );
  DFFQX1TS \Mem_reg[35][9]  ( .D(N1937), .CK(clk), .Q(\Mem[35][9] ) );
  DFFQX1TS \Mem_reg[35][8]  ( .D(N1936), .CK(clk), .Q(\Mem[35][8] ) );
  DFFQX1TS \Mem_reg[35][7]  ( .D(N1935), .CK(clk), .Q(\Mem[35][7] ) );
  DFFQX1TS \Mem_reg[35][6]  ( .D(N1934), .CK(clk), .Q(\Mem[35][6] ) );
  DFFQX1TS \Mem_reg[35][5]  ( .D(N1933), .CK(clk), .Q(\Mem[35][5] ) );
  DFFQX1TS \Mem_reg[35][4]  ( .D(N1932), .CK(clk), .Q(\Mem[35][4] ) );
  DFFQX1TS \Mem_reg[35][3]  ( .D(N1931), .CK(clk), .Q(\Mem[35][3] ) );
  DFFQX1TS \Mem_reg[35][2]  ( .D(N1930), .CK(clk), .Q(\Mem[35][2] ) );
  DFFQX1TS \Mem_reg[35][1]  ( .D(N1929), .CK(clk), .Q(\Mem[35][1] ) );
  DFFQX1TS \Mem_reg[35][0]  ( .D(N1928), .CK(clk), .Q(\Mem[35][0] ) );
  TLATXLTS \data_outA_reg[29]  ( .G(N162), .D(N63), .Q(data_outA[29]) );
  TLATXLTS \data_outA_reg[19]  ( .G(N162), .D(N73), .Q(data_outA[19]) );
  TLATXLTS \data_outA_reg[16]  ( .G(N162), .D(n520), .Q(data_outA[16]) );
  TLATXLTS \data_outA_reg[14]  ( .G(RAA[5]), .D(n519), .Q(data_outA[14]) );
  TLATXLTS \data_outA_reg[9]  ( .G(N162), .D(N83), .Q(data_outA[9]) );
  TLATXLTS \data_outA_reg[4]  ( .G(N162), .D(n514), .Q(data_outA[4]) );
  TLATXLTS \data_outA_reg[8]  ( .G(N162), .D(n516), .Q(data_outA[8]) );
  TLATXLTS \data_outA_reg[26]  ( .G(N162), .D(N66), .Q(data_outA[26]) );
  TLATXLTS \data_outA_reg[25]  ( .G(N162), .D(N67), .Q(data_outA[25]) );
  TLATXLTS \data_outA_reg[23]  ( .G(N162), .D(N69), .Q(data_outA[23]) );
  TLATXLTS \data_outA_reg[31]  ( .G(N162), .D(n525), .Q(data_outA[31]) );
  TLATXLTS \data_outA_reg[30]  ( .G(RAA[5]), .D(n524), .Q(data_outA[30]) );
  TLATXLTS \data_outA_reg[28]  ( .G(N162), .D(N64), .Q(data_outA[28]) );
  TLATXLTS \data_outA_reg[27]  ( .G(RAA[5]), .D(N65), .Q(data_outA[27]) );
  TLATXLTS \data_outA_reg[20]  ( .G(RAA[5]), .D(n522), .Q(data_outA[20]) );
  TLATXLTS \data_outA_reg[22]  ( .G(N162), .D(n523), .Q(data_outA[22]) );
  TLATXLTS \data_outA_reg[21]  ( .G(N162), .D(N71), .Q(data_outA[21]) );
  TLATXLTS \data_outA_reg[18]  ( .G(RAA[5]), .D(n521), .Q(data_outA[18]) );
  TLATXLTS \data_outA_reg[17]  ( .G(RAA[5]), .D(N75), .Q(data_outA[17]) );
  TLATXLTS \data_outA_reg[15]  ( .G(N162), .D(N77), .Q(data_outA[15]) );
  TLATXLTS \data_outA_reg[13]  ( .G(RAA[5]), .D(N79), .Q(data_outA[13]) );
  TLATXLTS \data_outA_reg[12]  ( .G(N162), .D(n518), .Q(data_outA[12]) );
  TLATXLTS \data_outA_reg[11]  ( .G(N162), .D(N81), .Q(data_outA[11]) );
  TLATXLTS \data_outA_reg[10]  ( .G(RAA[5]), .D(n517), .Q(data_outA[10]) );
  TLATXLTS \data_outA_reg[7]  ( .G(RAA[5]), .D(N85), .Q(data_outA[7]) );
  TLATXLTS \data_outA_reg[6]  ( .G(N162), .D(n515), .Q(data_outA[6]) );
  TLATXLTS \data_outA_reg[5]  ( .G(N162), .D(N87), .Q(data_outA[5]) );
  TLATXLTS \data_outA_reg[1]  ( .G(N162), .D(N91), .Q(data_outA[1]) );
  TLATXLTS \data_outA_reg[0]  ( .G(N162), .D(N92), .Q(data_outA[0]) );
  TLATXLTS \data_outA_reg[3]  ( .G(N162), .D(N89), .Q(data_outA[3]) );
  TLATXLTS \data_outA_reg[2]  ( .G(N162), .D(n513), .Q(data_outA[2]) );
  TLATXLTS \data_outA_reg[24]  ( .G(N162), .D(N68), .Q(data_outA[24]) );
  DFFQX1TS \Mem_reg[33][31]  ( .D(n407), .CK(clk), .Q(\Mem[33][31] ) );
  DFFQX1TS \Mem_reg[33][30]  ( .D(n406), .CK(clk), .Q(\Mem[33][30] ) );
  DFFQX1TS \Mem_reg[33][29]  ( .D(n405), .CK(clk), .Q(\Mem[33][29] ) );
  DFFQX1TS \Mem_reg[33][28]  ( .D(n404), .CK(clk), .Q(\Mem[33][28] ) );
  DFFQX1TS \Mem_reg[33][27]  ( .D(n403), .CK(clk), .Q(\Mem[33][27] ) );
  DFFQX1TS \Mem_reg[33][26]  ( .D(n402), .CK(clk), .Q(\Mem[33][26] ) );
  DFFQX1TS \Mem_reg[33][25]  ( .D(n401), .CK(clk), .Q(\Mem[33][25] ) );
  DFFQX1TS \Mem_reg[33][24]  ( .D(n400), .CK(clk), .Q(\Mem[33][24] ) );
  DFFQX1TS \Mem_reg[33][23]  ( .D(n399), .CK(clk), .Q(\Mem[33][23] ) );
  DFFQX1TS \Mem_reg[33][22]  ( .D(n398), .CK(clk), .Q(\Mem[33][22] ) );
  DFFQX1TS \Mem_reg[33][21]  ( .D(n397), .CK(clk), .Q(\Mem[33][21] ) );
  DFFQX1TS \Mem_reg[33][20]  ( .D(n396), .CK(clk), .Q(\Mem[33][20] ) );
  DFFQX1TS \Mem_reg[33][19]  ( .D(n395), .CK(clk), .Q(\Mem[33][19] ) );
  DFFQX1TS \Mem_reg[33][18]  ( .D(n394), .CK(clk), .Q(\Mem[33][18] ) );
  DFFQX1TS \Mem_reg[33][17]  ( .D(n393), .CK(clk), .Q(\Mem[33][17] ) );
  DFFQX1TS \Mem_reg[33][16]  ( .D(n392), .CK(clk), .Q(\Mem[33][16] ) );
  DFFQX1TS \Mem_reg[33][15]  ( .D(n391), .CK(clk), .Q(\Mem[33][15] ) );
  DFFQX1TS \Mem_reg[33][14]  ( .D(n390), .CK(clk), .Q(\Mem[33][14] ) );
  DFFQX1TS \Mem_reg[33][13]  ( .D(n389), .CK(clk), .Q(\Mem[33][13] ) );
  DFFQX1TS \Mem_reg[33][12]  ( .D(n388), .CK(clk), .Q(\Mem[33][12] ) );
  DFFQX1TS \Mem_reg[33][11]  ( .D(n387), .CK(clk), .Q(\Mem[33][11] ) );
  DFFQX1TS \Mem_reg[33][10]  ( .D(n386), .CK(clk), .Q(\Mem[33][10] ) );
  DFFQX1TS \Mem_reg[33][9]  ( .D(n385), .CK(clk), .Q(\Mem[33][9] ) );
  DFFQX1TS \Mem_reg[33][8]  ( .D(n384), .CK(clk), .Q(\Mem[33][8] ) );
  DFFQX1TS \Mem_reg[33][7]  ( .D(n383), .CK(clk), .Q(\Mem[33][7] ) );
  DFFQX1TS \Mem_reg[33][6]  ( .D(n382), .CK(clk), .Q(\Mem[33][6] ) );
  DFFQX1TS \Mem_reg[33][5]  ( .D(n381), .CK(clk), .Q(\Mem[33][5] ) );
  DFFQX1TS \Mem_reg[33][4]  ( .D(n380), .CK(clk), .Q(\Mem[33][4] ) );
  DFFQX1TS \Mem_reg[33][3]  ( .D(n379), .CK(clk), .Q(\Mem[33][3] ) );
  DFFQX1TS \Mem_reg[33][2]  ( .D(n378), .CK(clk), .Q(\Mem[33][2] ) );
  DFFQX1TS \Mem_reg[33][1]  ( .D(n377), .CK(clk), .Q(\Mem[33][1] ) );
  DFFQX1TS \Mem_reg[33][0]  ( .D(n376), .CK(clk), .Q(\Mem[33][0] ) );
  DFFQX1TS \Mem_reg[34][31]  ( .D(n439), .CK(clk), .Q(\Mem[34][31] ) );
  DFFQX1TS \Mem_reg[34][30]  ( .D(n438), .CK(clk), .Q(\Mem[34][30] ) );
  DFFQX1TS \Mem_reg[34][29]  ( .D(n437), .CK(clk), .Q(\Mem[34][29] ) );
  DFFQX1TS \Mem_reg[34][28]  ( .D(n436), .CK(clk), .Q(\Mem[34][28] ) );
  DFFQX1TS \Mem_reg[34][27]  ( .D(n435), .CK(clk), .Q(\Mem[34][27] ) );
  DFFQX1TS \Mem_reg[34][26]  ( .D(n434), .CK(clk), .Q(\Mem[34][26] ) );
  DFFQX1TS \Mem_reg[34][25]  ( .D(n433), .CK(clk), .Q(\Mem[34][25] ) );
  DFFQX1TS \Mem_reg[34][24]  ( .D(n432), .CK(clk), .Q(\Mem[34][24] ) );
  DFFQX1TS \Mem_reg[34][23]  ( .D(n431), .CK(clk), .Q(\Mem[34][23] ) );
  DFFQX1TS \Mem_reg[34][22]  ( .D(n430), .CK(clk), .Q(\Mem[34][22] ) );
  DFFQX1TS \Mem_reg[34][21]  ( .D(n429), .CK(clk), .Q(\Mem[34][21] ) );
  DFFQX1TS \Mem_reg[34][20]  ( .D(n428), .CK(clk), .Q(\Mem[34][20] ) );
  DFFQX1TS \Mem_reg[34][19]  ( .D(n427), .CK(clk), .Q(\Mem[34][19] ) );
  DFFQX1TS \Mem_reg[34][18]  ( .D(n426), .CK(clk), .Q(\Mem[34][18] ) );
  DFFQX1TS \Mem_reg[34][17]  ( .D(n425), .CK(clk), .Q(\Mem[34][17] ) );
  DFFQX1TS \Mem_reg[34][16]  ( .D(n424), .CK(clk), .Q(\Mem[34][16] ) );
  DFFQX1TS \Mem_reg[34][15]  ( .D(n423), .CK(clk), .Q(\Mem[34][15] ) );
  DFFQX1TS \Mem_reg[34][14]  ( .D(n422), .CK(clk), .Q(\Mem[34][14] ) );
  DFFQX1TS \Mem_reg[34][13]  ( .D(n421), .CK(clk), .Q(\Mem[34][13] ) );
  DFFQX1TS \Mem_reg[34][12]  ( .D(n420), .CK(clk), .Q(\Mem[34][12] ) );
  DFFQX1TS \Mem_reg[34][11]  ( .D(n419), .CK(clk), .Q(\Mem[34][11] ) );
  DFFQX1TS \Mem_reg[34][10]  ( .D(n418), .CK(clk), .Q(\Mem[34][10] ) );
  DFFQX1TS \Mem_reg[34][9]  ( .D(n417), .CK(clk), .Q(\Mem[34][9] ) );
  DFFQX1TS \Mem_reg[34][8]  ( .D(n416), .CK(clk), .Q(\Mem[34][8] ) );
  DFFQX1TS \Mem_reg[34][7]  ( .D(n415), .CK(clk), .Q(\Mem[34][7] ) );
  DFFQX1TS \Mem_reg[34][6]  ( .D(n414), .CK(clk), .Q(\Mem[34][6] ) );
  DFFQX1TS \Mem_reg[34][5]  ( .D(n413), .CK(clk), .Q(\Mem[34][5] ) );
  DFFQX1TS \Mem_reg[34][4]  ( .D(n412), .CK(clk), .Q(\Mem[34][4] ) );
  DFFQX1TS \Mem_reg[34][3]  ( .D(n411), .CK(clk), .Q(\Mem[34][3] ) );
  DFFQX1TS \Mem_reg[34][2]  ( .D(n410), .CK(clk), .Q(\Mem[34][2] ) );
  DFFQX1TS \Mem_reg[34][1]  ( .D(n409), .CK(clk), .Q(\Mem[34][1] ) );
  DFFQX1TS \Mem_reg[34][0]  ( .D(n408), .CK(clk), .Q(\Mem[34][0] ) );
  DFFQX1TS \Mem_reg[32][31]  ( .D(n375), .CK(clk), .Q(\Mem[32][31] ) );
  DFFQX1TS \Mem_reg[32][30]  ( .D(n374), .CK(clk), .Q(\Mem[32][30] ) );
  DFFQX1TS \Mem_reg[32][29]  ( .D(n373), .CK(clk), .Q(\Mem[32][29] ) );
  DFFQX1TS \Mem_reg[32][28]  ( .D(n372), .CK(clk), .Q(\Mem[32][28] ) );
  DFFQX1TS \Mem_reg[32][27]  ( .D(n371), .CK(clk), .Q(\Mem[32][27] ) );
  DFFQX1TS \Mem_reg[32][26]  ( .D(n370), .CK(clk), .Q(\Mem[32][26] ) );
  DFFQX1TS \Mem_reg[32][25]  ( .D(n369), .CK(clk), .Q(\Mem[32][25] ) );
  DFFQX1TS \Mem_reg[32][24]  ( .D(n368), .CK(clk), .Q(\Mem[32][24] ) );
  DFFQX1TS \Mem_reg[32][23]  ( .D(n367), .CK(clk), .Q(\Mem[32][23] ) );
  DFFQX1TS \Mem_reg[32][22]  ( .D(n366), .CK(clk), .Q(\Mem[32][22] ) );
  DFFQX1TS \Mem_reg[32][21]  ( .D(n365), .CK(clk), .Q(\Mem[32][21] ) );
  DFFQX1TS \Mem_reg[32][20]  ( .D(n364), .CK(clk), .Q(\Mem[32][20] ) );
  DFFQX1TS \Mem_reg[32][19]  ( .D(n363), .CK(clk), .Q(\Mem[32][19] ) );
  DFFQX1TS \Mem_reg[32][18]  ( .D(n362), .CK(clk), .Q(\Mem[32][18] ) );
  DFFQX1TS \Mem_reg[32][17]  ( .D(n361), .CK(clk), .Q(\Mem[32][17] ) );
  DFFQX1TS \Mem_reg[32][16]  ( .D(n360), .CK(clk), .Q(\Mem[32][16] ) );
  DFFQX1TS \Mem_reg[32][15]  ( .D(n359), .CK(clk), .Q(\Mem[32][15] ) );
  DFFQX1TS \Mem_reg[32][14]  ( .D(n358), .CK(clk), .Q(\Mem[32][14] ) );
  DFFQX1TS \Mem_reg[32][13]  ( .D(n357), .CK(clk), .Q(\Mem[32][13] ) );
  DFFQX1TS \Mem_reg[32][12]  ( .D(n356), .CK(clk), .Q(\Mem[32][12] ) );
  DFFQX1TS \Mem_reg[32][11]  ( .D(n355), .CK(clk), .Q(\Mem[32][11] ) );
  DFFQX1TS \Mem_reg[32][10]  ( .D(n354), .CK(clk), .Q(\Mem[32][10] ) );
  DFFQX1TS \Mem_reg[32][9]  ( .D(n353), .CK(clk), .Q(\Mem[32][9] ) );
  DFFQX1TS \Mem_reg[32][8]  ( .D(n352), .CK(clk), .Q(\Mem[32][8] ) );
  DFFQX1TS \Mem_reg[32][7]  ( .D(n351), .CK(clk), .Q(\Mem[32][7] ) );
  DFFQX1TS \Mem_reg[32][6]  ( .D(n350), .CK(clk), .Q(\Mem[32][6] ) );
  DFFQX1TS \Mem_reg[32][5]  ( .D(n349), .CK(clk), .Q(\Mem[32][5] ) );
  DFFQX1TS \Mem_reg[32][4]  ( .D(n348), .CK(clk), .Q(\Mem[32][4] ) );
  DFFQX1TS \Mem_reg[32][3]  ( .D(n347), .CK(clk), .Q(\Mem[32][3] ) );
  DFFQX1TS \Mem_reg[32][2]  ( .D(n346), .CK(clk), .Q(\Mem[32][2] ) );
  DFFQX1TS \Mem_reg[32][1]  ( .D(n345), .CK(clk), .Q(\Mem[32][1] ) );
  DFFQX1TS \Mem_reg[32][0]  ( .D(n344), .CK(clk), .Q(\Mem[32][0] ) );
  NOR2X4TS U3 ( .A(n130), .B(n4), .Y(n444) );
  NOR2X4TS U4 ( .A(n132), .B(n4), .Y(n456) );
  NOR2X4TS U5 ( .A(n135), .B(n4), .Y(n443) );
  NOR2X4TS U6 ( .A(n137), .B(n4), .Y(n455) );
  CLKAND2X2TS U7 ( .A(n70), .B(n44), .Y(n45) );
  NAND3X2TS U8 ( .A(WA[0]), .B(WA[5]), .C(n477), .Y(n476) );
  NAND3BX2TS U9 ( .AN(WA[0]), .B(WA[5]), .C(WA[1]), .Y(n475) );
  NAND3BX2TS U10 ( .AN(WA[0]), .B(WA[5]), .C(n477), .Y(n478) );
  NAND2BX2TS U11 ( .AN(enable[1]), .B(N162), .Y(n526) );
  NOR2X4TS U12 ( .A(n39), .B(n11), .Y(n105) );
  NOR2X4TS U13 ( .A(n38), .B(n11), .Y(n106) );
  NOR2X4TS U14 ( .A(n43), .B(n11), .Y(n107) );
  NOR2X4TS U15 ( .A(n42), .B(n11), .Y(n108) );
  INVX2TS U16 ( .A(data_in[31]), .Y(n479) );
  NAND3X1TS U17 ( .A(WA[1]), .B(WA[0]), .C(WA[5]), .Y(n473) );
  NOR2XLTS U18 ( .A(n479), .B(n473), .Y(N1959) );
  INVX2TS U19 ( .A(data_in[15]), .Y(n495) );
  NOR2XLTS U20 ( .A(n495), .B(n473), .Y(N1943) );
  INVX2TS U21 ( .A(data_in[0]), .Y(n510) );
  NOR2XLTS U22 ( .A(n510), .B(n473), .Y(N1928) );
  INVX2TS U23 ( .A(data_in[22]), .Y(n488) );
  NOR2XLTS U24 ( .A(n488), .B(n473), .Y(N1950) );
  INVX2TS U25 ( .A(data_in[5]), .Y(n505) );
  NOR2XLTS U26 ( .A(n505), .B(n473), .Y(N1933) );
  INVX2TS U27 ( .A(data_in[21]), .Y(n489) );
  NOR2XLTS U28 ( .A(n489), .B(n473), .Y(N1949) );
  INVX2TS U29 ( .A(data_in[18]), .Y(n492) );
  NOR2XLTS U30 ( .A(n492), .B(n473), .Y(N1946) );
  INVX2TS U31 ( .A(data_in[6]), .Y(n504) );
  NOR2XLTS U32 ( .A(n504), .B(n473), .Y(N1934) );
  INVX2TS U33 ( .A(data_in[13]), .Y(n497) );
  NOR2XLTS U34 ( .A(n497), .B(n473), .Y(N1941) );
  INVX2TS U35 ( .A(data_in[19]), .Y(n491) );
  NOR2XLTS U36 ( .A(n491), .B(n473), .Y(N1947) );
  INVX2TS U37 ( .A(data_in[9]), .Y(n501) );
  NOR2XLTS U38 ( .A(n501), .B(n473), .Y(N1937) );
  INVX2TS U39 ( .A(data_in[4]), .Y(n506) );
  NOR2XLTS U40 ( .A(n506), .B(n473), .Y(N1932) );
  INVX2TS U41 ( .A(data_in[24]), .Y(n486) );
  NOR2XLTS U42 ( .A(n486), .B(n473), .Y(N1952) );
  INVX2TS U43 ( .A(data_in[23]), .Y(n487) );
  NOR2XLTS U44 ( .A(n487), .B(n473), .Y(N1951) );
  INVX2TS U45 ( .A(data_in[25]), .Y(n485) );
  NOR2XLTS U46 ( .A(n485), .B(n473), .Y(N1953) );
  INVX2TS U47 ( .A(data_in[26]), .Y(n484) );
  NOR2XLTS U48 ( .A(n484), .B(n473), .Y(N1954) );
  INVX2TS U49 ( .A(data_in[27]), .Y(n483) );
  NOR2XLTS U50 ( .A(n483), .B(n473), .Y(N1955) );
  INVX2TS U51 ( .A(data_in[28]), .Y(n482) );
  NOR2XLTS U52 ( .A(n482), .B(n473), .Y(N1956) );
  INVX2TS U53 ( .A(data_in[29]), .Y(n481) );
  NOR2XLTS U54 ( .A(n481), .B(n473), .Y(N1957) );
  INVX2TS U55 ( .A(RAB[0]), .Y(n3) );
  INVX2TS U56 ( .A(RAB[1]), .Y(n2) );
  NAND2X1TS U57 ( .A(n3), .B(n2), .Y(n135) );
  NOR2BX1TS U58 ( .AN(RAB[5]), .B(RAB[4]), .Y(n1) );
  NOR2XLTS U59 ( .A(RAB[2]), .B(RAB[3]), .Y(n114) );
  NAND2X1TS U60 ( .A(n1), .B(n114), .Y(n4) );
  NAND2X1TS U61 ( .A(RAB[0]), .B(n2), .Y(n137) );
  AOI22X1TS U62 ( .A0(n443), .A1(\Mem[32][30] ), .B0(n455), .B1(\Mem[33][30] ), 
        .Y(n6) );
  NAND2X1TS U63 ( .A(RAB[1]), .B(n3), .Y(n130) );
  NAND2X1TS U64 ( .A(RAB[0]), .B(RAB[1]), .Y(n132) );
  AOI22X1TS U65 ( .A0(n444), .A1(\Mem[34][30] ), .B0(n456), .B1(\Mem[35][30] ), 
        .Y(n5) );
  NAND2X1TS U66 ( .A(n6), .B(n5), .Y(n511) );
  AOI22X1TS U67 ( .A0(n443), .A1(\Mem[32][31] ), .B0(n455), .B1(\Mem[33][31] ), 
        .Y(n8) );
  AOI22X1TS U68 ( .A0(n444), .A1(\Mem[34][31] ), .B0(n456), .B1(\Mem[35][31] ), 
        .Y(n7) );
  NAND2X1TS U69 ( .A(n8), .B(n7), .Y(n512) );
  INVX2TS U70 ( .A(RAA[0]), .Y(n10) );
  INVX2TS U71 ( .A(RAA[1]), .Y(n9) );
  NAND2X1TS U72 ( .A(n10), .B(n9), .Y(n38) );
  INVX2TS U73 ( .A(RAA[5]), .Y(n11) );
  NAND2X1TS U74 ( .A(RAA[0]), .B(n9), .Y(n39) );
  AOI22X1TS U75 ( .A0(n106), .A1(\Mem[32][2] ), .B0(n105), .B1(\Mem[33][2] ), 
        .Y(n13) );
  NAND2X1TS U76 ( .A(RAA[1]), .B(n10), .Y(n42) );
  NAND2X1TS U77 ( .A(RAA[0]), .B(RAA[1]), .Y(n43) );
  AOI22X1TS U78 ( .A0(n108), .A1(\Mem[34][2] ), .B0(n107), .B1(\Mem[35][2] ), 
        .Y(n12) );
  NAND2X1TS U79 ( .A(n13), .B(n12), .Y(n513) );
  AOI22X1TS U80 ( .A0(n106), .A1(\Mem[32][4] ), .B0(n105), .B1(\Mem[33][4] ), 
        .Y(n15) );
  AOI22X1TS U81 ( .A0(n108), .A1(\Mem[34][4] ), .B0(n107), .B1(\Mem[35][4] ), 
        .Y(n14) );
  NAND2X1TS U82 ( .A(n15), .B(n14), .Y(n514) );
  AOI22X1TS U83 ( .A0(n106), .A1(\Mem[32][6] ), .B0(n105), .B1(\Mem[33][6] ), 
        .Y(n17) );
  AOI22X1TS U84 ( .A0(n108), .A1(\Mem[34][6] ), .B0(n107), .B1(\Mem[35][6] ), 
        .Y(n16) );
  NAND2X1TS U85 ( .A(n17), .B(n16), .Y(n515) );
  AOI22X1TS U86 ( .A0(n106), .A1(\Mem[32][8] ), .B0(n105), .B1(\Mem[33][8] ), 
        .Y(n19) );
  AOI22X1TS U87 ( .A0(n108), .A1(\Mem[34][8] ), .B0(n107), .B1(\Mem[35][8] ), 
        .Y(n18) );
  NAND2X1TS U88 ( .A(n19), .B(n18), .Y(n516) );
  AOI22X1TS U89 ( .A0(n106), .A1(\Mem[32][10] ), .B0(n105), .B1(\Mem[33][10] ), 
        .Y(n21) );
  AOI22X1TS U90 ( .A0(n108), .A1(\Mem[34][10] ), .B0(n107), .B1(\Mem[35][10] ), 
        .Y(n20) );
  NAND2X1TS U91 ( .A(n21), .B(n20), .Y(n517) );
  AOI22X1TS U92 ( .A0(n106), .A1(\Mem[32][12] ), .B0(n105), .B1(\Mem[33][12] ), 
        .Y(n23) );
  AOI22X1TS U93 ( .A0(n108), .A1(\Mem[34][12] ), .B0(n107), .B1(\Mem[35][12] ), 
        .Y(n22) );
  NAND2X1TS U94 ( .A(n23), .B(n22), .Y(n518) );
  AOI22X1TS U95 ( .A0(n106), .A1(\Mem[32][14] ), .B0(n105), .B1(\Mem[33][14] ), 
        .Y(n25) );
  AOI22X1TS U96 ( .A0(n108), .A1(\Mem[34][14] ), .B0(n107), .B1(\Mem[35][14] ), 
        .Y(n24) );
  NAND2X1TS U97 ( .A(n25), .B(n24), .Y(n519) );
  AOI22X1TS U98 ( .A0(n106), .A1(\Mem[32][16] ), .B0(n105), .B1(\Mem[33][16] ), 
        .Y(n27) );
  AOI22X1TS U99 ( .A0(n108), .A1(\Mem[34][16] ), .B0(n107), .B1(\Mem[35][16] ), 
        .Y(n26) );
  NAND2X1TS U100 ( .A(n27), .B(n26), .Y(n520) );
  AOI22X1TS U101 ( .A0(n106), .A1(\Mem[32][18] ), .B0(n105), .B1(\Mem[33][18] ), .Y(n29) );
  AOI22X1TS U102 ( .A0(n108), .A1(\Mem[34][18] ), .B0(n107), .B1(\Mem[35][18] ), .Y(n28) );
  NAND2X1TS U103 ( .A(n29), .B(n28), .Y(n521) );
  AOI22X1TS U104 ( .A0(n106), .A1(\Mem[32][20] ), .B0(n105), .B1(\Mem[33][20] ), .Y(n31) );
  AOI22X1TS U105 ( .A0(n108), .A1(\Mem[34][20] ), .B0(n107), .B1(\Mem[35][20] ), .Y(n30) );
  NAND2X1TS U106 ( .A(n31), .B(n30), .Y(n522) );
  AOI22X1TS U107 ( .A0(n106), .A1(\Mem[32][22] ), .B0(n105), .B1(\Mem[33][22] ), .Y(n33) );
  AOI22X1TS U108 ( .A0(n108), .A1(\Mem[34][22] ), .B0(n107), .B1(\Mem[35][22] ), .Y(n32) );
  NAND2X1TS U109 ( .A(n33), .B(n32), .Y(n523) );
  AOI22X1TS U110 ( .A0(n106), .A1(\Mem[32][30] ), .B0(n105), .B1(\Mem[33][30] ), .Y(n35) );
  AOI22X1TS U111 ( .A0(n108), .A1(\Mem[34][30] ), .B0(n107), .B1(\Mem[35][30] ), .Y(n34) );
  NAND2X1TS U112 ( .A(n35), .B(n34), .Y(n524) );
  AOI22X1TS U113 ( .A0(n106), .A1(\Mem[32][31] ), .B0(n105), .B1(\Mem[33][31] ), .Y(n37) );
  AOI22X1TS U114 ( .A0(n108), .A1(\Mem[34][31] ), .B0(n107), .B1(\Mem[35][31] ), .Y(n36) );
  NAND2X1TS U115 ( .A(n37), .B(n36), .Y(n525) );
  NOR2XLTS U116 ( .A(n38), .B(RAA[5]), .Y(n41) );
  NOR2XLTS U117 ( .A(n39), .B(RAA[5]), .Y(n40) );
  NOR2XLTS U118 ( .A(n41), .B(n40), .Y(n70) );
  NOR2XLTS U119 ( .A(n42), .B(RAA[5]), .Y(n61) );
  NOR2XLTS U120 ( .A(n43), .B(RAA[5]), .Y(n71) );
  NOR2XLTS U121 ( .A(n61), .B(n71), .Y(n44) );
  AOI22X1TS U122 ( .A0(n106), .A1(\Mem[32][29] ), .B0(n105), .B1(\Mem[33][29] ), .Y(n47) );
  AOI22X1TS U123 ( .A0(n108), .A1(\Mem[34][29] ), .B0(n107), .B1(\Mem[35][29] ), .Y(n46) );
  CLKAND2X2TS U124 ( .A(n47), .B(n46), .Y(n48) );
  NAND2X1TS U125 ( .A(n45), .B(n48), .Y(N63) );
  AOI22X1TS U126 ( .A0(n106), .A1(\Mem[32][28] ), .B0(n105), .B1(\Mem[33][28] ), .Y(n50) );
  AOI22X1TS U127 ( .A0(n108), .A1(\Mem[34][28] ), .B0(n107), .B1(\Mem[35][28] ), .Y(n49) );
  CLKAND2X2TS U128 ( .A(n50), .B(n49), .Y(n51) );
  NAND2X1TS U129 ( .A(n45), .B(n51), .Y(N64) );
  AOI22X1TS U130 ( .A0(n106), .A1(\Mem[32][27] ), .B0(n105), .B1(\Mem[33][27] ), .Y(n53) );
  AOI22X1TS U131 ( .A0(n108), .A1(\Mem[34][27] ), .B0(n107), .B1(\Mem[35][27] ), .Y(n52) );
  CLKAND2X2TS U132 ( .A(n53), .B(n52), .Y(n54) );
  NAND2X1TS U133 ( .A(n45), .B(n54), .Y(N65) );
  AOI22X1TS U134 ( .A0(n106), .A1(\Mem[32][26] ), .B0(n105), .B1(\Mem[33][26] ), .Y(n56) );
  AOI22X1TS U135 ( .A0(n108), .A1(\Mem[34][26] ), .B0(n107), .B1(\Mem[35][26] ), .Y(n55) );
  CLKAND2X2TS U136 ( .A(n56), .B(n55), .Y(n57) );
  NAND2X1TS U137 ( .A(n45), .B(n57), .Y(N66) );
  AOI22X1TS U138 ( .A0(n106), .A1(\Mem[32][25] ), .B0(n105), .B1(\Mem[33][25] ), .Y(n59) );
  AOI22X1TS U139 ( .A0(n108), .A1(\Mem[34][25] ), .B0(n107), .B1(\Mem[35][25] ), .Y(n58) );
  CLKAND2X2TS U140 ( .A(n59), .B(n58), .Y(n60) );
  NAND2X1TS U141 ( .A(n45), .B(n60), .Y(N67) );
  INVX2TS U142 ( .A(n61), .Y(n62) );
  CLKAND2X2TS U143 ( .A(n70), .B(n62), .Y(n66) );
  AOI22X1TS U144 ( .A0(n106), .A1(\Mem[32][24] ), .B0(n105), .B1(\Mem[33][24] ), .Y(n64) );
  AOI22X1TS U145 ( .A0(n108), .A1(\Mem[34][24] ), .B0(n107), .B1(\Mem[35][24] ), .Y(n63) );
  CLKAND2X2TS U146 ( .A(n64), .B(n63), .Y(n65) );
  NAND2X1TS U147 ( .A(n66), .B(n65), .Y(N68) );
  AOI22X1TS U148 ( .A0(n106), .A1(\Mem[32][23] ), .B0(n105), .B1(\Mem[33][23] ), .Y(n68) );
  AOI22X1TS U149 ( .A0(n108), .A1(\Mem[34][23] ), .B0(n107), .B1(\Mem[35][23] ), .Y(n67) );
  CLKAND2X2TS U150 ( .A(n68), .B(n67), .Y(n69) );
  NAND2X1TS U151 ( .A(n70), .B(n69), .Y(N69) );
  INVX2TS U152 ( .A(n71), .Y(n112) );
  AOI22X1TS U153 ( .A0(n106), .A1(\Mem[32][21] ), .B0(n105), .B1(\Mem[33][21] ), .Y(n73) );
  AOI22X1TS U154 ( .A0(n108), .A1(\Mem[34][21] ), .B0(n107), .B1(\Mem[35][21] ), .Y(n72) );
  CLKAND2X2TS U155 ( .A(n73), .B(n72), .Y(n74) );
  NAND2X1TS U156 ( .A(n112), .B(n74), .Y(N71) );
  AOI22X1TS U157 ( .A0(n106), .A1(\Mem[32][19] ), .B0(n105), .B1(\Mem[33][19] ), .Y(n76) );
  AOI22X1TS U158 ( .A0(n108), .A1(\Mem[34][19] ), .B0(n107), .B1(\Mem[35][19] ), .Y(n75) );
  CLKAND2X2TS U159 ( .A(n76), .B(n75), .Y(n77) );
  NAND2X1TS U160 ( .A(n112), .B(n77), .Y(N73) );
  AOI22X1TS U161 ( .A0(n106), .A1(\Mem[32][17] ), .B0(n105), .B1(\Mem[33][17] ), .Y(n79) );
  AOI22X1TS U162 ( .A0(n108), .A1(\Mem[34][17] ), .B0(n107), .B1(\Mem[35][17] ), .Y(n78) );
  CLKAND2X2TS U163 ( .A(n79), .B(n78), .Y(n80) );
  NAND2X1TS U164 ( .A(n112), .B(n80), .Y(N75) );
  AOI22X1TS U165 ( .A0(n106), .A1(\Mem[32][15] ), .B0(n105), .B1(\Mem[33][15] ), .Y(n82) );
  AOI22X1TS U166 ( .A0(n108), .A1(\Mem[34][15] ), .B0(n107), .B1(\Mem[35][15] ), .Y(n81) );
  CLKAND2X2TS U167 ( .A(n82), .B(n81), .Y(n83) );
  NAND2X1TS U168 ( .A(n112), .B(n83), .Y(N77) );
  AOI22X1TS U169 ( .A0(n106), .A1(\Mem[32][13] ), .B0(n105), .B1(\Mem[33][13] ), .Y(n85) );
  AOI22X1TS U170 ( .A0(n108), .A1(\Mem[34][13] ), .B0(n107), .B1(\Mem[35][13] ), .Y(n84) );
  CLKAND2X2TS U171 ( .A(n85), .B(n84), .Y(n86) );
  NAND2X1TS U172 ( .A(n112), .B(n86), .Y(N79) );
  AOI22X1TS U173 ( .A0(n106), .A1(\Mem[32][11] ), .B0(n105), .B1(\Mem[33][11] ), .Y(n88) );
  AOI22X1TS U174 ( .A0(n108), .A1(\Mem[34][11] ), .B0(n107), .B1(\Mem[35][11] ), .Y(n87) );
  CLKAND2X2TS U175 ( .A(n88), .B(n87), .Y(n89) );
  NAND2X1TS U176 ( .A(n112), .B(n89), .Y(N81) );
  AOI22X1TS U177 ( .A0(n106), .A1(\Mem[32][9] ), .B0(n105), .B1(\Mem[33][9] ), 
        .Y(n91) );
  AOI22X1TS U178 ( .A0(n108), .A1(\Mem[34][9] ), .B0(n107), .B1(\Mem[35][9] ), 
        .Y(n90) );
  CLKAND2X2TS U179 ( .A(n91), .B(n90), .Y(n92) );
  NAND2X1TS U180 ( .A(n112), .B(n92), .Y(N83) );
  AOI22X1TS U181 ( .A0(n106), .A1(\Mem[32][7] ), .B0(n105), .B1(\Mem[33][7] ), 
        .Y(n94) );
  AOI22X1TS U182 ( .A0(n108), .A1(\Mem[34][7] ), .B0(n107), .B1(\Mem[35][7] ), 
        .Y(n93) );
  CLKAND2X2TS U183 ( .A(n94), .B(n93), .Y(n95) );
  NAND2X1TS U184 ( .A(n112), .B(n95), .Y(N85) );
  AOI22X1TS U185 ( .A0(n106), .A1(\Mem[32][5] ), .B0(n105), .B1(\Mem[33][5] ), 
        .Y(n97) );
  AOI22X1TS U186 ( .A0(n108), .A1(\Mem[34][5] ), .B0(n107), .B1(\Mem[35][5] ), 
        .Y(n96) );
  CLKAND2X2TS U187 ( .A(n97), .B(n96), .Y(n98) );
  NAND2X1TS U188 ( .A(n112), .B(n98), .Y(N87) );
  AOI22X1TS U189 ( .A0(n106), .A1(\Mem[32][3] ), .B0(n105), .B1(\Mem[33][3] ), 
        .Y(n100) );
  AOI22X1TS U190 ( .A0(n108), .A1(\Mem[34][3] ), .B0(n107), .B1(\Mem[35][3] ), 
        .Y(n99) );
  CLKAND2X2TS U191 ( .A(n100), .B(n99), .Y(n101) );
  NAND2X1TS U192 ( .A(n112), .B(n101), .Y(N89) );
  AOI22X1TS U193 ( .A0(n106), .A1(\Mem[32][1] ), .B0(n105), .B1(\Mem[33][1] ), 
        .Y(n103) );
  AOI22X1TS U194 ( .A0(n108), .A1(\Mem[34][1] ), .B0(n107), .B1(\Mem[35][1] ), 
        .Y(n102) );
  CLKAND2X2TS U195 ( .A(n103), .B(n102), .Y(n104) );
  NAND2X1TS U196 ( .A(n112), .B(n104), .Y(N91) );
  AOI22X1TS U197 ( .A0(n106), .A1(\Mem[32][0] ), .B0(n105), .B1(\Mem[33][0] ), 
        .Y(n110) );
  AOI22X1TS U198 ( .A0(n108), .A1(\Mem[34][0] ), .B0(n107), .B1(\Mem[35][0] ), 
        .Y(n109) );
  CLKAND2X2TS U199 ( .A(n110), .B(n109), .Y(n111) );
  NAND2X1TS U200 ( .A(n112), .B(n111), .Y(N92) );
  NOR2BX1TS U201 ( .AN(RAB[4]), .B(RAB[5]), .Y(n133) );
  NAND2X1TS U202 ( .A(n114), .B(n133), .Y(n113) );
  NOR2XLTS U203 ( .A(n130), .B(n113), .Y(n156) );
  NOR2XLTS U204 ( .A(n132), .B(n113), .Y(n168) );
  NOR2XLTS U205 ( .A(n156), .B(n168), .Y(n310) );
  NOR2BX1TS U206 ( .AN(RAB[2]), .B(RAB[3]), .Y(n118) );
  NAND2X1TS U207 ( .A(n118), .B(n133), .Y(n131) );
  NOR2XLTS U208 ( .A(n135), .B(n131), .Y(n191) );
  INVX2TS U209 ( .A(n191), .Y(n293) );
  NOR2XLTS U210 ( .A(n135), .B(n113), .Y(n144) );
  NOR2XLTS U211 ( .A(n137), .B(n113), .Y(n155) );
  NOR2X1TS U212 ( .A(n144), .B(n155), .Y(n335) );
  NAND3XLTS U213 ( .A(n310), .B(n293), .C(n335), .Y(n125) );
  NOR2XLTS U214 ( .A(RAB[4]), .B(RAB[5]), .Y(n122) );
  NAND2X1TS U215 ( .A(n114), .B(n122), .Y(n117) );
  NOR2XLTS U216 ( .A(n135), .B(n117), .Y(n115) );
  NOR2XLTS U217 ( .A(n137), .B(n117), .Y(n116) );
  NOR2XLTS U218 ( .A(n115), .B(n116), .Y(n189) );
  NOR2XLTS U219 ( .A(n130), .B(n117), .Y(n177) );
  NOR2XLTS U220 ( .A(n132), .B(n117), .Y(n205) );
  NOR2XLTS U221 ( .A(n177), .B(n205), .Y(n165) );
  NAND2X1TS U222 ( .A(n118), .B(n122), .Y(n120) );
  NOR2XLTS U223 ( .A(n135), .B(n120), .Y(n178) );
  NOR2XLTS U224 ( .A(n137), .B(n120), .Y(n119) );
  NOR2XLTS U225 ( .A(n178), .B(n119), .Y(n270) );
  NOR2XLTS U226 ( .A(n130), .B(n120), .Y(n313) );
  NOR2XLTS U227 ( .A(n132), .B(n120), .Y(n281) );
  NOR2XLTS U228 ( .A(n313), .B(n281), .Y(n269) );
  NAND4XLTS U229 ( .A(n189), .B(n165), .C(n270), .D(n269), .Y(n147) );
  NOR2BX1TS U230 ( .AN(RAB[3]), .B(RAB[2]), .Y(n134) );
  NAND2X1TS U231 ( .A(n134), .B(n122), .Y(n121) );
  NOR2XLTS U232 ( .A(n135), .B(n121), .Y(n181) );
  NOR2XLTS U233 ( .A(n137), .B(n121), .Y(n207) );
  NOR2X1TS U234 ( .A(n181), .B(n207), .Y(n464) );
  NOR2XLTS U235 ( .A(n130), .B(n121), .Y(n153) );
  NOR2XLTS U236 ( .A(n132), .B(n121), .Y(n166) );
  NOR2X1TS U237 ( .A(n153), .B(n166), .Y(n450) );
  NAND3XLTS U238 ( .A(RAB[2]), .B(RAB[3]), .C(n122), .Y(n123) );
  NOR2XLTS U239 ( .A(n135), .B(n123), .Y(n220) );
  NOR2XLTS U240 ( .A(n137), .B(n123), .Y(n145) );
  NOR2XLTS U241 ( .A(n220), .B(n145), .Y(n286) );
  NOR2XLTS U242 ( .A(n130), .B(n123), .Y(n154) );
  NOR2XLTS U243 ( .A(n132), .B(n123), .Y(n167) );
  NOR2X1TS U244 ( .A(n154), .B(n167), .Y(n461) );
  NAND4XLTS U245 ( .A(n464), .B(n450), .C(n286), .D(n461), .Y(n124) );
  NOR3XLTS U246 ( .A(n125), .B(n147), .C(n124), .Y(n129) );
  AOI22X1TS U247 ( .A0(n443), .A1(\Mem[32][29] ), .B0(n455), .B1(\Mem[33][29] ), .Y(n127) );
  AOI22X1TS U248 ( .A0(n444), .A1(\Mem[34][29] ), .B0(n456), .B1(\Mem[35][29] ), .Y(n126) );
  CLKAND2X2TS U249 ( .A(n127), .B(n126), .Y(n128) );
  NAND2X1TS U250 ( .A(n129), .B(n128), .Y(N95) );
  INVX2TS U251 ( .A(n220), .Y(n276) );
  NAND3XLTS U252 ( .A(n450), .B(n276), .C(n464), .Y(n139) );
  NOR2XLTS U253 ( .A(n137), .B(n131), .Y(n190) );
  INVX2TS U254 ( .A(n190), .Y(n278) );
  NOR2XLTS U255 ( .A(n130), .B(n131), .Y(n157) );
  NOR2XLTS U256 ( .A(n132), .B(n131), .Y(n169) );
  NOR2XLTS U257 ( .A(n157), .B(n169), .Y(n302) );
  NAND2X1TS U258 ( .A(n278), .B(n302), .Y(n138) );
  NAND2X1TS U259 ( .A(n134), .B(n133), .Y(n136) );
  NOR2XLTS U260 ( .A(n135), .B(n136), .Y(n303) );
  NOR2X1TS U261 ( .A(n137), .B(n136), .Y(n451) );
  OR2X1TS U262 ( .A(n303), .B(n451), .Y(n465) );
  NOR4XLTS U263 ( .A(n147), .B(n139), .C(n138), .D(n465), .Y(n143) );
  AOI22X1TS U264 ( .A0(n443), .A1(\Mem[32][28] ), .B0(n455), .B1(\Mem[33][28] ), .Y(n141) );
  AOI22X1TS U265 ( .A0(n444), .A1(\Mem[34][28] ), .B0(n456), .B1(\Mem[35][28] ), .Y(n140) );
  CLKAND2X2TS U266 ( .A(n141), .B(n140), .Y(n142) );
  NAND2X1TS U267 ( .A(n143), .B(n142), .Y(N96) );
  INVX2TS U268 ( .A(n144), .Y(n301) );
  NAND3XLTS U269 ( .A(n278), .B(n302), .C(n301), .Y(n148) );
  INVX2TS U270 ( .A(n145), .Y(n462) );
  NAND2X1TS U271 ( .A(n462), .B(n461), .Y(n146) );
  NOR3XLTS U272 ( .A(n148), .B(n147), .C(n146), .Y(n152) );
  AOI22X1TS U273 ( .A0(n443), .A1(\Mem[32][27] ), .B0(n455), .B1(\Mem[33][27] ), .Y(n150) );
  AOI22X1TS U274 ( .A0(n444), .A1(\Mem[34][27] ), .B0(n456), .B1(\Mem[35][27] ), .Y(n149) );
  CLKAND2X2TS U275 ( .A(n150), .B(n149), .Y(n151) );
  NAND2X1TS U276 ( .A(n152), .B(n151), .Y(N97) );
  NAND3XLTS U277 ( .A(n165), .B(n270), .C(n189), .Y(n160) );
  INVX2TS U278 ( .A(n153), .Y(n440) );
  INVX2TS U279 ( .A(n154), .Y(n318) );
  NAND4XLTS U280 ( .A(n464), .B(n440), .C(n462), .D(n318), .Y(n159) );
  INVX2TS U281 ( .A(n155), .Y(n243) );
  INVX2TS U282 ( .A(n156), .Y(n294) );
  INVX2TS U283 ( .A(n157), .Y(n332) );
  NAND4XLTS U284 ( .A(n243), .B(n294), .C(n278), .D(n332), .Y(n158) );
  NOR4XLTS U285 ( .A(n160), .B(n159), .C(n158), .D(n465), .Y(n164) );
  AOI22X1TS U286 ( .A0(n443), .A1(\Mem[32][26] ), .B0(n455), .B1(\Mem[33][26] ), .Y(n162) );
  AOI22X1TS U287 ( .A0(n444), .A1(\Mem[34][26] ), .B0(n456), .B1(\Mem[35][26] ), .Y(n161) );
  CLKAND2X2TS U288 ( .A(n162), .B(n161), .Y(n163) );
  NAND2X1TS U289 ( .A(n164), .B(n163), .Y(N98) );
  INVX2TS U290 ( .A(n313), .Y(n206) );
  NAND3XLTS U291 ( .A(n165), .B(n206), .C(n189), .Y(n172) );
  INVX2TS U292 ( .A(n166), .Y(n463) );
  INVX2TS U293 ( .A(n167), .Y(n449) );
  NAND4XLTS U294 ( .A(n464), .B(n463), .C(n462), .D(n449), .Y(n171) );
  INVX2TS U295 ( .A(n168), .Y(n334) );
  INVX2TS U296 ( .A(n169), .Y(n277) );
  NAND4XLTS U297 ( .A(n243), .B(n334), .C(n278), .D(n277), .Y(n170) );
  NOR4XLTS U298 ( .A(n172), .B(n171), .C(n170), .D(n303), .Y(n176) );
  AOI22X1TS U299 ( .A0(n443), .A1(\Mem[32][25] ), .B0(n455), .B1(\Mem[33][25] ), .Y(n174) );
  AOI22X1TS U300 ( .A0(n444), .A1(\Mem[34][25] ), .B0(n456), .B1(\Mem[35][25] ), .Y(n173) );
  CLKAND2X2TS U301 ( .A(n174), .B(n173), .Y(n175) );
  NAND2X1TS U302 ( .A(n176), .B(n175), .Y(N99) );
  INVX2TS U303 ( .A(n177), .Y(n180) );
  INVX2TS U304 ( .A(n178), .Y(n256) );
  INVX2TS U305 ( .A(n281), .Y(n179) );
  NAND4XLTS U306 ( .A(n189), .B(n180), .C(n256), .D(n179), .Y(n184) );
  INVX2TS U307 ( .A(n181), .Y(n199) );
  NAND3XLTS U308 ( .A(n286), .B(n461), .C(n199), .Y(n183) );
  NAND2X1TS U309 ( .A(n335), .B(n310), .Y(n182) );
  NOR4XLTS U310 ( .A(n184), .B(n183), .C(n182), .D(n465), .Y(n188) );
  AOI22X1TS U311 ( .A0(n443), .A1(\Mem[32][24] ), .B0(n455), .B1(\Mem[33][24] ), .Y(n186) );
  AOI22X1TS U312 ( .A0(n444), .A1(\Mem[34][24] ), .B0(n456), .B1(\Mem[35][24] ), .Y(n185) );
  CLKAND2X2TS U313 ( .A(n186), .B(n185), .Y(n187) );
  NAND2X1TS U314 ( .A(n188), .B(n187), .Y(N100) );
  NAND2X1TS U315 ( .A(n189), .B(n206), .Y(n194) );
  NAND2X1TS U316 ( .A(n199), .B(n450), .Y(n193) );
  NOR2XLTS U317 ( .A(n191), .B(n190), .Y(n333) );
  NAND2X1TS U318 ( .A(n333), .B(n332), .Y(n192) );
  NOR4XLTS U319 ( .A(n194), .B(n193), .C(n192), .D(n465), .Y(n198) );
  AOI22X1TS U320 ( .A0(n443), .A1(\Mem[32][23] ), .B0(n455), .B1(\Mem[33][23] ), .Y(n196) );
  AOI22X1TS U321 ( .A0(n444), .A1(\Mem[34][23] ), .B0(n456), .B1(\Mem[35][23] ), .Y(n195) );
  CLKAND2X2TS U322 ( .A(n196), .B(n195), .Y(n197) );
  NAND2X1TS U323 ( .A(n198), .B(n197), .Y(N101) );
  NAND3XLTS U324 ( .A(n463), .B(n461), .C(n199), .Y(n200) );
  NAND2X1TS U325 ( .A(n335), .B(n293), .Y(n441) );
  NOR4XLTS U326 ( .A(n281), .B(n200), .C(n441), .D(n303), .Y(n204) );
  AOI22X1TS U327 ( .A0(n443), .A1(\Mem[32][22] ), .B0(n455), .B1(\Mem[33][22] ), .Y(n202) );
  AOI22X1TS U328 ( .A0(n444), .A1(\Mem[34][22] ), .B0(n456), .B1(\Mem[35][22] ), .Y(n201) );
  CLKAND2X2TS U329 ( .A(n202), .B(n201), .Y(n203) );
  NAND2X1TS U330 ( .A(n204), .B(n203), .Y(N102) );
  INVX2TS U331 ( .A(n205), .Y(n268) );
  NAND3XLTS U332 ( .A(n256), .B(n206), .C(n268), .Y(n321) );
  INVX2TS U333 ( .A(n207), .Y(n343) );
  NAND2X1TS U334 ( .A(n343), .B(n462), .Y(n209) );
  NAND3XLTS U335 ( .A(n333), .B(n277), .C(n294), .Y(n208) );
  NOR4XLTS U336 ( .A(n321), .B(n209), .C(n208), .D(n303), .Y(n213) );
  AOI22X1TS U337 ( .A0(n443), .A1(\Mem[32][21] ), .B0(n455), .B1(\Mem[33][21] ), .Y(n211) );
  AOI22X1TS U338 ( .A0(n444), .A1(\Mem[34][21] ), .B0(n456), .B1(\Mem[35][21] ), .Y(n210) );
  CLKAND2X2TS U339 ( .A(n211), .B(n210), .Y(n212) );
  NAND2X1TS U340 ( .A(n213), .B(n212), .Y(N103) );
  INVX2TS U341 ( .A(n269), .Y(n296) );
  NAND4XLTS U342 ( .A(n464), .B(n450), .C(n462), .D(n449), .Y(n215) );
  NAND4XLTS U343 ( .A(n301), .B(n310), .C(n333), .D(n277), .Y(n214) );
  NOR4XLTS U344 ( .A(n296), .B(n215), .C(n214), .D(n465), .Y(n219) );
  AOI22X1TS U345 ( .A0(n443), .A1(\Mem[32][20] ), .B0(n455), .B1(\Mem[33][20] ), .Y(n217) );
  AOI22X1TS U346 ( .A0(n444), .A1(\Mem[34][20] ), .B0(n456), .B1(\Mem[35][20] ), .Y(n216) );
  CLKAND2X2TS U347 ( .A(n217), .B(n216), .Y(n218) );
  NAND2X1TS U348 ( .A(n219), .B(n218), .Y(N104) );
  NAND2X1TS U349 ( .A(n268), .B(n270), .Y(n337) );
  NAND3XLTS U350 ( .A(n276), .B(n318), .C(n343), .Y(n221) );
  NAND3XLTS U351 ( .A(n278), .B(n277), .C(n243), .Y(n319) );
  NOR4XLTS U352 ( .A(n337), .B(n221), .C(n319), .D(n465), .Y(n225) );
  AOI22X1TS U353 ( .A0(n443), .A1(\Mem[32][19] ), .B0(n455), .B1(\Mem[33][19] ), .Y(n223) );
  AOI22X1TS U354 ( .A0(n444), .A1(\Mem[34][19] ), .B0(n456), .B1(\Mem[35][19] ), .Y(n222) );
  CLKAND2X2TS U355 ( .A(n223), .B(n222), .Y(n224) );
  NAND2X1TS U356 ( .A(n225), .B(n224), .Y(N105) );
  NAND3XLTS U357 ( .A(n276), .B(n449), .C(n463), .Y(n226) );
  NAND3XLTS U358 ( .A(n310), .B(n332), .C(n301), .Y(n452) );
  NOR4XLTS U359 ( .A(n313), .B(n226), .C(n452), .D(n451), .Y(n230) );
  AOI22X1TS U360 ( .A0(n443), .A1(\Mem[32][18] ), .B0(n455), .B1(\Mem[33][18] ), .Y(n228) );
  AOI22X1TS U361 ( .A0(n444), .A1(\Mem[34][18] ), .B0(n456), .B1(\Mem[35][18] ), .Y(n227) );
  CLKAND2X2TS U362 ( .A(n228), .B(n227), .Y(n229) );
  NAND2X1TS U363 ( .A(n230), .B(n229), .Y(N106) );
  NAND3XLTS U364 ( .A(n276), .B(n449), .C(n450), .Y(n232) );
  NAND4XLTS U365 ( .A(n335), .B(n334), .C(n293), .D(n302), .Y(n231) );
  NOR4XLTS U366 ( .A(n321), .B(n232), .C(n231), .D(n451), .Y(n236) );
  AOI22X1TS U367 ( .A0(n443), .A1(\Mem[32][17] ), .B0(n455), .B1(\Mem[33][17] ), .Y(n234) );
  AOI22X1TS U368 ( .A0(n444), .A1(\Mem[34][17] ), .B0(n456), .B1(\Mem[35][17] ), .Y(n233) );
  CLKAND2X2TS U369 ( .A(n234), .B(n233), .Y(n235) );
  NAND2X1TS U370 ( .A(n236), .B(n235), .Y(N107) );
  NAND3XLTS U371 ( .A(n276), .B(n461), .C(n450), .Y(n238) );
  NAND3XLTS U372 ( .A(n334), .B(n277), .C(n301), .Y(n237) );
  NOR3XLTS U373 ( .A(n465), .B(n238), .C(n237), .Y(n242) );
  AOI22X1TS U374 ( .A0(n443), .A1(\Mem[32][16] ), .B0(n455), .B1(\Mem[33][16] ), .Y(n240) );
  AOI22X1TS U375 ( .A0(n444), .A1(\Mem[34][16] ), .B0(n456), .B1(\Mem[35][16] ), .Y(n239) );
  CLKAND2X2TS U376 ( .A(n240), .B(n239), .Y(n241) );
  NAND2X1TS U377 ( .A(n242), .B(n241), .Y(N108) );
  NAND4XLTS U378 ( .A(n343), .B(n440), .C(n462), .D(n318), .Y(n245) );
  NAND3XLTS U379 ( .A(n334), .B(n333), .C(n243), .Y(n244) );
  NOR4XLTS U380 ( .A(n337), .B(n245), .C(n244), .D(n451), .Y(n249) );
  AOI22X1TS U381 ( .A0(n443), .A1(\Mem[32][15] ), .B0(n455), .B1(\Mem[33][15] ), .Y(n247) );
  AOI22X1TS U382 ( .A0(n444), .A1(\Mem[34][15] ), .B0(n456), .B1(\Mem[35][15] ), .Y(n246) );
  CLKAND2X2TS U383 ( .A(n247), .B(n246), .Y(n248) );
  NAND2X1TS U384 ( .A(n249), .B(n248), .Y(N109) );
  NAND4XLTS U385 ( .A(n343), .B(n440), .C(n276), .D(n318), .Y(n251) );
  NAND2X1TS U386 ( .A(n278), .B(n332), .Y(n250) );
  NOR3XLTS U387 ( .A(n303), .B(n251), .C(n250), .Y(n255) );
  AOI22X1TS U388 ( .A0(n443), .A1(\Mem[32][14] ), .B0(n455), .B1(\Mem[33][14] ), .Y(n253) );
  AOI22X1TS U389 ( .A0(n444), .A1(\Mem[34][14] ), .B0(n456), .B1(\Mem[35][14] ), .Y(n252) );
  CLKAND2X2TS U390 ( .A(n253), .B(n252), .Y(n254) );
  NAND2X1TS U391 ( .A(n255), .B(n254), .Y(N110) );
  NAND2X1TS U392 ( .A(n268), .B(n256), .Y(n454) );
  NAND4XLTS U393 ( .A(n343), .B(n450), .C(n276), .D(n449), .Y(n336) );
  NAND4XLTS U394 ( .A(n301), .B(n334), .C(n293), .D(n332), .Y(n257) );
  NOR4XLTS U395 ( .A(n454), .B(n336), .C(n257), .D(n303), .Y(n261) );
  AOI22X1TS U396 ( .A0(n443), .A1(\Mem[32][13] ), .B0(n455), .B1(\Mem[33][13] ), .Y(n259) );
  AOI22X1TS U397 ( .A0(n444), .A1(\Mem[34][13] ), .B0(n456), .B1(\Mem[35][13] ), .Y(n258) );
  CLKAND2X2TS U398 ( .A(n259), .B(n258), .Y(n260) );
  NAND2X1TS U399 ( .A(n261), .B(n260), .Y(N111) );
  NAND3XLTS U400 ( .A(n286), .B(n449), .C(n450), .Y(n263) );
  NAND4XLTS U401 ( .A(n335), .B(n294), .C(n278), .D(n332), .Y(n262) );
  NOR3XLTS U402 ( .A(n451), .B(n263), .C(n262), .Y(n267) );
  AOI22X1TS U403 ( .A0(n443), .A1(\Mem[32][12] ), .B0(n455), .B1(\Mem[33][12] ), .Y(n265) );
  AOI22X1TS U404 ( .A0(n444), .A1(\Mem[34][12] ), .B0(n456), .B1(\Mem[35][12] ), .Y(n264) );
  CLKAND2X2TS U405 ( .A(n265), .B(n264), .Y(n266) );
  NAND2X1TS U406 ( .A(n267), .B(n266), .Y(N112) );
  NAND3XLTS U407 ( .A(n270), .B(n269), .C(n268), .Y(n468) );
  NAND2X1TS U408 ( .A(n464), .B(n461), .Y(n295) );
  NAND3XLTS U409 ( .A(n278), .B(n277), .C(n301), .Y(n271) );
  NOR4XLTS U410 ( .A(n468), .B(n295), .C(n271), .D(n451), .Y(n275) );
  AOI22X1TS U411 ( .A0(n443), .A1(\Mem[32][11] ), .B0(n455), .B1(\Mem[33][11] ), .Y(n273) );
  AOI22X1TS U412 ( .A0(n444), .A1(\Mem[34][11] ), .B0(n456), .B1(\Mem[35][11] ), .Y(n272) );
  CLKAND2X2TS U413 ( .A(n273), .B(n272), .Y(n274) );
  NAND2X1TS U414 ( .A(n275), .B(n274), .Y(N113) );
  NAND3XLTS U415 ( .A(n276), .B(n449), .C(n464), .Y(n280) );
  NAND4XLTS U416 ( .A(n335), .B(n334), .C(n278), .D(n277), .Y(n279) );
  NOR4XLTS U417 ( .A(n281), .B(n280), .C(n279), .D(n465), .Y(n285) );
  AOI22X1TS U418 ( .A0(n443), .A1(\Mem[32][10] ), .B0(n455), .B1(\Mem[33][10] ), .Y(n283) );
  AOI22X1TS U419 ( .A0(n444), .A1(\Mem[34][10] ), .B0(n456), .B1(\Mem[35][10] ), .Y(n282) );
  CLKAND2X2TS U420 ( .A(n283), .B(n282), .Y(n284) );
  NAND2X1TS U421 ( .A(n285), .B(n284), .Y(N114) );
  NAND4XLTS U422 ( .A(n343), .B(n450), .C(n286), .D(n461), .Y(n288) );
  NAND2X1TS U423 ( .A(n335), .B(n294), .Y(n287) );
  NOR4XLTS U424 ( .A(n321), .B(n288), .C(n287), .D(n465), .Y(n292) );
  AOI22X1TS U425 ( .A0(n443), .A1(\Mem[32][9] ), .B0(n455), .B1(\Mem[33][9] ), 
        .Y(n290) );
  AOI22X1TS U426 ( .A0(n444), .A1(\Mem[34][9] ), .B0(n456), .B1(\Mem[35][9] ), 
        .Y(n289) );
  CLKAND2X2TS U427 ( .A(n290), .B(n289), .Y(n291) );
  NAND2X1TS U428 ( .A(n292), .B(n291), .Y(N115) );
  NAND4XLTS U429 ( .A(n301), .B(n294), .C(n293), .D(n302), .Y(n466) );
  NOR4XLTS U430 ( .A(n296), .B(n295), .C(n466), .D(n303), .Y(n300) );
  AOI22X1TS U431 ( .A0(n443), .A1(\Mem[32][8] ), .B0(n455), .B1(\Mem[33][8] ), 
        .Y(n298) );
  AOI22X1TS U432 ( .A0(n444), .A1(\Mem[34][8] ), .B0(n456), .B1(\Mem[35][8] ), 
        .Y(n297) );
  CLKAND2X2TS U433 ( .A(n298), .B(n297), .Y(n299) );
  NAND2X1TS U434 ( .A(n300), .B(n299), .Y(N116) );
  NAND3XLTS U435 ( .A(n276), .B(n461), .C(n343), .Y(n305) );
  NAND3XLTS U436 ( .A(n310), .B(n302), .C(n301), .Y(n304) );
  NOR4XLTS U437 ( .A(n337), .B(n305), .C(n304), .D(n303), .Y(n309) );
  AOI22X1TS U438 ( .A0(n443), .A1(\Mem[32][7] ), .B0(n455), .B1(\Mem[33][7] ), 
        .Y(n307) );
  AOI22X1TS U439 ( .A0(n444), .A1(\Mem[34][7] ), .B0(n456), .B1(\Mem[35][7] ), 
        .Y(n306) );
  CLKAND2X2TS U440 ( .A(n307), .B(n306), .Y(n308) );
  NAND2X1TS U441 ( .A(n309), .B(n308), .Y(N117) );
  NAND3XLTS U442 ( .A(n440), .B(n276), .C(n343), .Y(n312) );
  NAND3XLTS U443 ( .A(n333), .B(n332), .C(n310), .Y(n311) );
  NOR4XLTS U444 ( .A(n313), .B(n312), .C(n311), .D(n451), .Y(n317) );
  AOI22X1TS U445 ( .A0(n443), .A1(\Mem[32][6] ), .B0(n455), .B1(\Mem[33][6] ), 
        .Y(n315) );
  AOI22X1TS U446 ( .A0(n444), .A1(\Mem[34][6] ), .B0(n456), .B1(\Mem[35][6] ), 
        .Y(n314) );
  CLKAND2X2TS U447 ( .A(n315), .B(n314), .Y(n316) );
  NAND2X1TS U448 ( .A(n317), .B(n316), .Y(N118) );
  NAND4XLTS U449 ( .A(n343), .B(n450), .C(n462), .D(n318), .Y(n320) );
  NOR4XLTS U450 ( .A(n321), .B(n320), .C(n319), .D(n451), .Y(n325) );
  AOI22X1TS U451 ( .A0(n443), .A1(\Mem[32][5] ), .B0(n455), .B1(\Mem[33][5] ), 
        .Y(n323) );
  AOI22X1TS U452 ( .A0(n444), .A1(\Mem[34][5] ), .B0(n456), .B1(\Mem[35][5] ), 
        .Y(n322) );
  CLKAND2X2TS U453 ( .A(n323), .B(n322), .Y(n324) );
  NAND2X1TS U454 ( .A(n325), .B(n324), .Y(N119) );
  NAND3XLTS U455 ( .A(n334), .B(n333), .C(n335), .Y(n327) );
  NAND3XLTS U456 ( .A(n462), .B(n449), .C(n440), .Y(n326) );
  NOR2XLTS U457 ( .A(n327), .B(n326), .Y(n331) );
  AOI22X1TS U458 ( .A0(n443), .A1(\Mem[32][4] ), .B0(n455), .B1(\Mem[33][4] ), 
        .Y(n329) );
  AOI22X1TS U459 ( .A0(n444), .A1(\Mem[34][4] ), .B0(n456), .B1(\Mem[35][4] ), 
        .Y(n328) );
  CLKAND2X2TS U460 ( .A(n329), .B(n328), .Y(n330) );
  NAND2X1TS U461 ( .A(n331), .B(n330), .Y(N120) );
  NAND4XLTS U462 ( .A(n335), .B(n334), .C(n333), .D(n332), .Y(n338) );
  NOR3XLTS U463 ( .A(n338), .B(n337), .C(n336), .Y(n342) );
  AOI22X1TS U464 ( .A0(n443), .A1(\Mem[32][3] ), .B0(n455), .B1(\Mem[33][3] ), 
        .Y(n340) );
  AOI22X1TS U465 ( .A0(n444), .A1(\Mem[34][3] ), .B0(n456), .B1(\Mem[35][3] ), 
        .Y(n339) );
  CLKAND2X2TS U466 ( .A(n340), .B(n339), .Y(n341) );
  NAND2X1TS U467 ( .A(n342), .B(n341), .Y(N121) );
  NAND3XLTS U468 ( .A(n440), .B(n461), .C(n343), .Y(n442) );
  NOR3XLTS U469 ( .A(n451), .B(n442), .C(n441), .Y(n448) );
  AOI22X1TS U470 ( .A0(n443), .A1(\Mem[32][2] ), .B0(n455), .B1(\Mem[33][2] ), 
        .Y(n446) );
  AOI22X1TS U471 ( .A0(n444), .A1(\Mem[34][2] ), .B0(n456), .B1(\Mem[35][2] ), 
        .Y(n445) );
  CLKAND2X2TS U472 ( .A(n446), .B(n445), .Y(n447) );
  NAND2X1TS U473 ( .A(n448), .B(n447), .Y(N122) );
  NAND2X1TS U474 ( .A(n450), .B(n449), .Y(n453) );
  NOR4XLTS U475 ( .A(n454), .B(n453), .C(n452), .D(n451), .Y(n460) );
  AOI22X1TS U476 ( .A0(n443), .A1(\Mem[32][1] ), .B0(n455), .B1(\Mem[33][1] ), 
        .Y(n458) );
  AOI22X1TS U477 ( .A0(n444), .A1(\Mem[34][1] ), .B0(n456), .B1(\Mem[35][1] ), 
        .Y(n457) );
  CLKAND2X2TS U478 ( .A(n458), .B(n457), .Y(n459) );
  NAND2X1TS U479 ( .A(n460), .B(n459), .Y(N123) );
  NAND4XLTS U480 ( .A(n464), .B(n463), .C(n462), .D(n461), .Y(n467) );
  NOR4XLTS U481 ( .A(n468), .B(n467), .C(n466), .D(n465), .Y(n472) );
  AOI22X1TS U482 ( .A0(n443), .A1(\Mem[32][0] ), .B0(n455), .B1(\Mem[33][0] ), 
        .Y(n470) );
  AOI22X1TS U483 ( .A0(n444), .A1(\Mem[34][0] ), .B0(n456), .B1(\Mem[35][0] ), 
        .Y(n469) );
  CLKAND2X2TS U484 ( .A(n470), .B(n469), .Y(n471) );
  NAND2X1TS U485 ( .A(n472), .B(n471), .Y(N124) );
  INVX2TS U486 ( .A(n473), .Y(n474) );
  INVX2TS U487 ( .A(data_in[1]), .Y(n509) );
  NAND2X1TS U488 ( .A(n474), .B(n509), .Y(N1929) );
  INVX2TS U489 ( .A(data_in[2]), .Y(n508) );
  NAND2X1TS U490 ( .A(n474), .B(n508), .Y(N1930) );
  INVX2TS U491 ( .A(data_in[3]), .Y(n507) );
  NAND2X1TS U492 ( .A(n474), .B(n507), .Y(N1931) );
  INVX2TS U493 ( .A(data_in[7]), .Y(n503) );
  NAND2X1TS U494 ( .A(n474), .B(n503), .Y(N1935) );
  INVX2TS U495 ( .A(data_in[8]), .Y(n502) );
  NAND2X1TS U496 ( .A(n474), .B(n502), .Y(N1936) );
  INVX2TS U497 ( .A(data_in[10]), .Y(n500) );
  NAND2X1TS U498 ( .A(n474), .B(n500), .Y(N1938) );
  INVX2TS U499 ( .A(data_in[11]), .Y(n499) );
  NAND2X1TS U500 ( .A(n474), .B(n499), .Y(N1939) );
  INVX2TS U501 ( .A(data_in[12]), .Y(n498) );
  NAND2X1TS U502 ( .A(n474), .B(n498), .Y(N1940) );
  INVX2TS U503 ( .A(data_in[14]), .Y(n496) );
  NAND2X1TS U504 ( .A(n474), .B(n496), .Y(N1942) );
  INVX2TS U505 ( .A(data_in[16]), .Y(n494) );
  NAND2X1TS U506 ( .A(n474), .B(n494), .Y(N1944) );
  INVX2TS U507 ( .A(data_in[17]), .Y(n493) );
  NAND2X1TS U508 ( .A(n474), .B(n493), .Y(N1945) );
  INVX2TS U509 ( .A(data_in[20]), .Y(n490) );
  NAND2X1TS U510 ( .A(n474), .B(n490), .Y(N1948) );
  INVX2TS U511 ( .A(data_in[30]), .Y(n480) );
  NAND2X1TS U512 ( .A(n474), .B(n480), .Y(N1958) );
  OAI2BB2XLTS U513 ( .B0(n475), .B1(n479), .A0N(n475), .A1N(\Mem[34][31] ), 
        .Y(n439) );
  OAI2BB2XLTS U514 ( .B0(n475), .B1(n480), .A0N(n475), .A1N(\Mem[34][30] ), 
        .Y(n438) );
  OAI2BB2XLTS U515 ( .B0(n475), .B1(n481), .A0N(n475), .A1N(\Mem[34][29] ), 
        .Y(n437) );
  OAI2BB2XLTS U516 ( .B0(n475), .B1(n482), .A0N(n475), .A1N(\Mem[34][28] ), 
        .Y(n436) );
  OAI2BB2XLTS U517 ( .B0(n475), .B1(n483), .A0N(n475), .A1N(\Mem[34][27] ), 
        .Y(n435) );
  OAI2BB2XLTS U518 ( .B0(n475), .B1(n484), .A0N(n475), .A1N(\Mem[34][26] ), 
        .Y(n434) );
  OAI2BB2XLTS U519 ( .B0(n475), .B1(n485), .A0N(n475), .A1N(\Mem[34][25] ), 
        .Y(n433) );
  OAI2BB2XLTS U520 ( .B0(n475), .B1(n486), .A0N(n475), .A1N(\Mem[34][24] ), 
        .Y(n432) );
  OAI2BB2XLTS U521 ( .B0(n475), .B1(n487), .A0N(n475), .A1N(\Mem[34][23] ), 
        .Y(n431) );
  OAI2BB2XLTS U522 ( .B0(n475), .B1(n488), .A0N(n475), .A1N(\Mem[34][22] ), 
        .Y(n430) );
  OAI2BB2XLTS U523 ( .B0(n475), .B1(n489), .A0N(n475), .A1N(\Mem[34][21] ), 
        .Y(n429) );
  OAI2BB2XLTS U524 ( .B0(n475), .B1(n490), .A0N(n475), .A1N(\Mem[34][20] ), 
        .Y(n428) );
  OAI2BB2XLTS U525 ( .B0(n475), .B1(n491), .A0N(n475), .A1N(\Mem[34][19] ), 
        .Y(n427) );
  OAI2BB2XLTS U526 ( .B0(n475), .B1(n492), .A0N(n475), .A1N(\Mem[34][18] ), 
        .Y(n426) );
  OAI2BB2XLTS U527 ( .B0(n475), .B1(n493), .A0N(n475), .A1N(\Mem[34][17] ), 
        .Y(n425) );
  OAI2BB2XLTS U528 ( .B0(n475), .B1(n494), .A0N(n475), .A1N(\Mem[34][16] ), 
        .Y(n424) );
  OAI2BB2XLTS U529 ( .B0(n475), .B1(n495), .A0N(n475), .A1N(\Mem[34][15] ), 
        .Y(n423) );
  OAI2BB2XLTS U530 ( .B0(n475), .B1(n496), .A0N(n475), .A1N(\Mem[34][14] ), 
        .Y(n422) );
  OAI2BB2XLTS U531 ( .B0(n475), .B1(n497), .A0N(n475), .A1N(\Mem[34][13] ), 
        .Y(n421) );
  OAI2BB2XLTS U532 ( .B0(n475), .B1(n498), .A0N(n475), .A1N(\Mem[34][12] ), 
        .Y(n420) );
  OAI2BB2XLTS U533 ( .B0(n475), .B1(n499), .A0N(n475), .A1N(\Mem[34][11] ), 
        .Y(n419) );
  OAI2BB2XLTS U534 ( .B0(n475), .B1(n500), .A0N(n475), .A1N(\Mem[34][10] ), 
        .Y(n418) );
  OAI2BB2XLTS U535 ( .B0(n475), .B1(n501), .A0N(n475), .A1N(\Mem[34][9] ), .Y(
        n417) );
  OAI2BB2XLTS U536 ( .B0(n475), .B1(n502), .A0N(n475), .A1N(\Mem[34][8] ), .Y(
        n416) );
  OAI2BB2XLTS U537 ( .B0(n475), .B1(n503), .A0N(n475), .A1N(\Mem[34][7] ), .Y(
        n415) );
  OAI2BB2XLTS U538 ( .B0(n475), .B1(n504), .A0N(n475), .A1N(\Mem[34][6] ), .Y(
        n414) );
  OAI2BB2XLTS U539 ( .B0(n475), .B1(n505), .A0N(n475), .A1N(\Mem[34][5] ), .Y(
        n413) );
  OAI2BB2XLTS U540 ( .B0(n475), .B1(n506), .A0N(n475), .A1N(\Mem[34][4] ), .Y(
        n412) );
  OAI2BB2XLTS U541 ( .B0(n475), .B1(n507), .A0N(n475), .A1N(\Mem[34][3] ), .Y(
        n411) );
  OAI2BB2XLTS U542 ( .B0(n475), .B1(n508), .A0N(n475), .A1N(\Mem[34][2] ), .Y(
        n410) );
  OAI2BB2XLTS U543 ( .B0(n475), .B1(n509), .A0N(n475), .A1N(\Mem[34][1] ), .Y(
        n409) );
  OAI2BB2XLTS U544 ( .B0(n475), .B1(n510), .A0N(n475), .A1N(\Mem[34][0] ), .Y(
        n408) );
  INVX2TS U545 ( .A(WA[1]), .Y(n477) );
  OAI2BB2XLTS U546 ( .B0(n476), .B1(n479), .A0N(n476), .A1N(\Mem[33][31] ), 
        .Y(n407) );
  OAI2BB2XLTS U547 ( .B0(n476), .B1(n480), .A0N(n476), .A1N(\Mem[33][30] ), 
        .Y(n406) );
  OAI2BB2XLTS U548 ( .B0(n476), .B1(n481), .A0N(n476), .A1N(\Mem[33][29] ), 
        .Y(n405) );
  OAI2BB2XLTS U549 ( .B0(n476), .B1(n482), .A0N(n476), .A1N(\Mem[33][28] ), 
        .Y(n404) );
  OAI2BB2XLTS U550 ( .B0(n476), .B1(n483), .A0N(n476), .A1N(\Mem[33][27] ), 
        .Y(n403) );
  OAI2BB2XLTS U551 ( .B0(n476), .B1(n484), .A0N(n476), .A1N(\Mem[33][26] ), 
        .Y(n402) );
  OAI2BB2XLTS U552 ( .B0(n476), .B1(n485), .A0N(n476), .A1N(\Mem[33][25] ), 
        .Y(n401) );
  OAI2BB2XLTS U553 ( .B0(n476), .B1(n486), .A0N(n476), .A1N(\Mem[33][24] ), 
        .Y(n400) );
  OAI2BB2XLTS U554 ( .B0(n476), .B1(n487), .A0N(n476), .A1N(\Mem[33][23] ), 
        .Y(n399) );
  OAI2BB2XLTS U555 ( .B0(n476), .B1(n488), .A0N(n476), .A1N(\Mem[33][22] ), 
        .Y(n398) );
  OAI2BB2XLTS U556 ( .B0(n476), .B1(n489), .A0N(n476), .A1N(\Mem[33][21] ), 
        .Y(n397) );
  OAI2BB2XLTS U557 ( .B0(n476), .B1(n490), .A0N(n476), .A1N(\Mem[33][20] ), 
        .Y(n396) );
  OAI2BB2XLTS U558 ( .B0(n476), .B1(n491), .A0N(n476), .A1N(\Mem[33][19] ), 
        .Y(n395) );
  OAI2BB2XLTS U559 ( .B0(n476), .B1(n492), .A0N(n476), .A1N(\Mem[33][18] ), 
        .Y(n394) );
  OAI2BB2XLTS U560 ( .B0(n476), .B1(n493), .A0N(n476), .A1N(\Mem[33][17] ), 
        .Y(n393) );
  OAI2BB2XLTS U561 ( .B0(n476), .B1(n494), .A0N(n476), .A1N(\Mem[33][16] ), 
        .Y(n392) );
  OAI2BB2XLTS U562 ( .B0(n476), .B1(n495), .A0N(n476), .A1N(\Mem[33][15] ), 
        .Y(n391) );
  OAI2BB2XLTS U563 ( .B0(n476), .B1(n496), .A0N(n476), .A1N(\Mem[33][14] ), 
        .Y(n390) );
  OAI2BB2XLTS U564 ( .B0(n476), .B1(n497), .A0N(n476), .A1N(\Mem[33][13] ), 
        .Y(n389) );
  OAI2BB2XLTS U565 ( .B0(n476), .B1(n498), .A0N(n476), .A1N(\Mem[33][12] ), 
        .Y(n388) );
  OAI2BB2XLTS U566 ( .B0(n476), .B1(n499), .A0N(n476), .A1N(\Mem[33][11] ), 
        .Y(n387) );
  OAI2BB2XLTS U567 ( .B0(n476), .B1(n500), .A0N(n476), .A1N(\Mem[33][10] ), 
        .Y(n386) );
  OAI2BB2XLTS U568 ( .B0(n476), .B1(n501), .A0N(n476), .A1N(\Mem[33][9] ), .Y(
        n385) );
  OAI2BB2XLTS U569 ( .B0(n476), .B1(n502), .A0N(n476), .A1N(\Mem[33][8] ), .Y(
        n384) );
  OAI2BB2XLTS U570 ( .B0(n476), .B1(n503), .A0N(n476), .A1N(\Mem[33][7] ), .Y(
        n383) );
  OAI2BB2XLTS U571 ( .B0(n476), .B1(n504), .A0N(n476), .A1N(\Mem[33][6] ), .Y(
        n382) );
  OAI2BB2XLTS U572 ( .B0(n476), .B1(n505), .A0N(n476), .A1N(\Mem[33][5] ), .Y(
        n381) );
  OAI2BB2XLTS U573 ( .B0(n476), .B1(n506), .A0N(n476), .A1N(\Mem[33][4] ), .Y(
        n380) );
  OAI2BB2XLTS U574 ( .B0(n476), .B1(n507), .A0N(n476), .A1N(\Mem[33][3] ), .Y(
        n379) );
  OAI2BB2XLTS U575 ( .B0(n476), .B1(n508), .A0N(n476), .A1N(\Mem[33][2] ), .Y(
        n378) );
  OAI2BB2XLTS U576 ( .B0(n476), .B1(n509), .A0N(n476), .A1N(\Mem[33][1] ), .Y(
        n377) );
  OAI2BB2XLTS U577 ( .B0(n476), .B1(n510), .A0N(n476), .A1N(\Mem[33][0] ), .Y(
        n376) );
  OAI2BB2XLTS U578 ( .B0(n478), .B1(n479), .A0N(n478), .A1N(\Mem[32][31] ), 
        .Y(n375) );
  OAI2BB2XLTS U579 ( .B0(n478), .B1(n480), .A0N(n478), .A1N(\Mem[32][30] ), 
        .Y(n374) );
  OAI2BB2XLTS U580 ( .B0(n478), .B1(n481), .A0N(n478), .A1N(\Mem[32][29] ), 
        .Y(n373) );
  OAI2BB2XLTS U581 ( .B0(n478), .B1(n482), .A0N(n478), .A1N(\Mem[32][28] ), 
        .Y(n372) );
  OAI2BB2XLTS U582 ( .B0(n478), .B1(n483), .A0N(n478), .A1N(\Mem[32][27] ), 
        .Y(n371) );
  OAI2BB2XLTS U583 ( .B0(n478), .B1(n484), .A0N(n478), .A1N(\Mem[32][26] ), 
        .Y(n370) );
  OAI2BB2XLTS U584 ( .B0(n478), .B1(n485), .A0N(n478), .A1N(\Mem[32][25] ), 
        .Y(n369) );
  OAI2BB2XLTS U585 ( .B0(n478), .B1(n486), .A0N(n478), .A1N(\Mem[32][24] ), 
        .Y(n368) );
  OAI2BB2XLTS U586 ( .B0(n478), .B1(n487), .A0N(n478), .A1N(\Mem[32][23] ), 
        .Y(n367) );
  OAI2BB2XLTS U587 ( .B0(n478), .B1(n488), .A0N(n478), .A1N(\Mem[32][22] ), 
        .Y(n366) );
  OAI2BB2XLTS U588 ( .B0(n478), .B1(n489), .A0N(n478), .A1N(\Mem[32][21] ), 
        .Y(n365) );
  OAI2BB2XLTS U589 ( .B0(n478), .B1(n490), .A0N(n478), .A1N(\Mem[32][20] ), 
        .Y(n364) );
  OAI2BB2XLTS U590 ( .B0(n478), .B1(n491), .A0N(n478), .A1N(\Mem[32][19] ), 
        .Y(n363) );
  OAI2BB2XLTS U591 ( .B0(n478), .B1(n492), .A0N(n478), .A1N(\Mem[32][18] ), 
        .Y(n362) );
  OAI2BB2XLTS U592 ( .B0(n478), .B1(n493), .A0N(n478), .A1N(\Mem[32][17] ), 
        .Y(n361) );
  OAI2BB2XLTS U593 ( .B0(n478), .B1(n494), .A0N(n478), .A1N(\Mem[32][16] ), 
        .Y(n360) );
  OAI2BB2XLTS U594 ( .B0(n478), .B1(n495), .A0N(n478), .A1N(\Mem[32][15] ), 
        .Y(n359) );
  OAI2BB2XLTS U595 ( .B0(n478), .B1(n496), .A0N(n478), .A1N(\Mem[32][14] ), 
        .Y(n358) );
  OAI2BB2XLTS U596 ( .B0(n478), .B1(n497), .A0N(n478), .A1N(\Mem[32][13] ), 
        .Y(n357) );
  OAI2BB2XLTS U597 ( .B0(n478), .B1(n498), .A0N(n478), .A1N(\Mem[32][12] ), 
        .Y(n356) );
  OAI2BB2XLTS U598 ( .B0(n478), .B1(n499), .A0N(n478), .A1N(\Mem[32][11] ), 
        .Y(n355) );
  OAI2BB2XLTS U599 ( .B0(n478), .B1(n500), .A0N(n478), .A1N(\Mem[32][10] ), 
        .Y(n354) );
  OAI2BB2XLTS U600 ( .B0(n478), .B1(n501), .A0N(n478), .A1N(\Mem[32][9] ), .Y(
        n353) );
  OAI2BB2XLTS U601 ( .B0(n478), .B1(n502), .A0N(n478), .A1N(\Mem[32][8] ), .Y(
        n352) );
  OAI2BB2XLTS U602 ( .B0(n478), .B1(n503), .A0N(n478), .A1N(\Mem[32][7] ), .Y(
        n351) );
  OAI2BB2XLTS U603 ( .B0(n478), .B1(n504), .A0N(n478), .A1N(\Mem[32][6] ), .Y(
        n350) );
  OAI2BB2XLTS U604 ( .B0(n478), .B1(n505), .A0N(n478), .A1N(\Mem[32][5] ), .Y(
        n349) );
  OAI2BB2XLTS U605 ( .B0(n478), .B1(n506), .A0N(n478), .A1N(\Mem[32][4] ), .Y(
        n348) );
  OAI2BB2XLTS U606 ( .B0(n478), .B1(n507), .A0N(n478), .A1N(\Mem[32][3] ), .Y(
        n347) );
  OAI2BB2XLTS U607 ( .B0(n478), .B1(n508), .A0N(n478), .A1N(\Mem[32][2] ), .Y(
        n346) );
  OAI2BB2XLTS U608 ( .B0(n478), .B1(n509), .A0N(n478), .A1N(\Mem[32][1] ), .Y(
        n345) );
  OAI2BB2XLTS U609 ( .B0(n478), .B1(n510), .A0N(n478), .A1N(\Mem[32][0] ), .Y(
        n344) );
endmodule


module FSM ( clk, reset, start, mq47, mp47, r31, msb, ms0_24, ms0_23, ms0_63, 
        comp1_g, comp2_g, stxor, st, sumor, mode, mux5, mux7, mux10, mux11, 
        mux15, mux16, mux18, mux19, mux22, mux23, mux1, mux4, mux6, mux12, 
        mux14, mux20, mux21, mux2, mux3, mux8, mux9, mux13, mux17, rf_we, 
        rf_rea, rf_reb, rf_wa, rf_raa, rf_rab, reg_sum, reg_i, reg_currterm, 
        reg_index, reg_reg, reg_r, reg_numbit, reg_e, reg_acc, reg_sc, reg_ec, 
        reg_mc, reg_sb, reg_eb, reg_mb, reg_sa, reg_ea, reg_ma, reg_sq, reg_eq, 
        reg_ss, reg_es, reg_ms, reg_st, reg_et, reg_sp, reg_ep, reg_es0, 
        reg_ss0, sr_res, sr_mq, sr_mt, sr_mp, ssr_ms0, alu1, alu2, counterii, 
        state );
  input [2:0] mode;
  output [1:0] mux1;
  output [1:0] mux4;
  output [1:0] mux6;
  output [1:0] mux12;
  output [1:0] mux14;
  output [1:0] mux20;
  output [1:0] mux21;
  output [2:0] mux2;
  output [2:0] mux3;
  output [2:0] mux8;
  output [2:0] mux9;
  output [2:0] mux13;
  output [2:0] mux17;
  output [5:0] rf_wa;
  output [5:0] rf_raa;
  output [5:0] rf_rab;
  output [1:0] sr_res;
  output [1:0] sr_mq;
  output [1:0] sr_mt;
  output [1:0] sr_mp;
  output [2:0] ssr_ms0;
  output [2:0] alu1;
  output [2:0] alu2;
  output [2:0] counterii;
  output [8:0] state;
  input clk, reset, start, mq47, mp47, r31, msb, ms0_24, ms0_23, ms0_63,
         comp1_g, comp2_g, stxor, st, sumor;
  output mux5, mux7, mux10, mux11, mux15, mux16, mux18, mux19, mux22, mux23,
         rf_we, rf_rea, rf_reb, reg_sum, reg_i, reg_currterm, reg_index,
         reg_reg, reg_r, reg_numbit, reg_e, reg_acc, reg_sc, reg_ec, reg_mc,
         reg_sb, reg_eb, reg_mb, reg_sa, reg_ea, reg_ma, reg_sq, reg_eq,
         reg_ss, reg_es, reg_ms, reg_st, reg_et, reg_sp, reg_ep, reg_es0,
         reg_ss0;
  wire   mux17_0, rf_wa_5, rf_rab_5, N2131, N2139, N2152, N2444, N2445, N2446,
         N2447, N2448, N2449, N2450, N2451, N2452, N2453, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660;
  wire   [8:0] nextstate;
  assign mux17[0] = mux17_0;
  assign rf_wa[5] = rf_wa_5;
  assign rf_rab[5] = rf_rab_5;
  assign N2131 = stxor;
  assign N2139 = mp47;
  assign N2152 = ms0_63;

  TLATXLTS \nextstate_reg[0]  ( .G(n660), .D(N2445), .Q(nextstate[0]) );
  TLATXLTS \nextstate_reg[7]  ( .G(n660), .D(N2452), .Q(nextstate[7]) );
  TLATXLTS \nextstate_reg[4]  ( .G(n660), .D(N2449), .Q(nextstate[4]) );
  TLATXLTS \nextstate_reg[6]  ( .G(n660), .D(N2451), .Q(nextstate[6]) );
  TLATXLTS \nextstate_reg[5]  ( .G(N2444), .D(N2450), .Q(nextstate[5]) );
  TLATXLTS \nextstate_reg[3]  ( .G(N2444), .D(N2448), .Q(nextstate[3]) );
  TLATXLTS \nextstate_reg[1]  ( .G(N2444), .D(N2446), .Q(nextstate[1]) );
  TLATXLTS \nextstate_reg[2]  ( .G(N2444), .D(N2447), .Q(nextstate[2]) );
  TLATXLTS \nextstate_reg[8]  ( .G(N2444), .D(N2453), .Q(nextstate[8]) );
  DFFQX1TS \state_reg[0]  ( .D(nextstate[0]), .CK(clk), .Q(state[0]) );
  DFFQX1TS \state_reg[1]  ( .D(nextstate[1]), .CK(clk), .Q(state[1]) );
  DFFQX1TS \state_reg[2]  ( .D(nextstate[2]), .CK(clk), .Q(state[2]) );
  DFFQX1TS \state_reg[4]  ( .D(nextstate[4]), .CK(clk), .Q(state[4]) );
  DFFQX1TS \state_reg[7]  ( .D(nextstate[7]), .CK(clk), .Q(state[7]) );
  DFFQX1TS \state_reg[5]  ( .D(nextstate[5]), .CK(clk), .Q(state[5]) );
  DFFQX1TS \state_reg[8]  ( .D(nextstate[8]), .CK(clk), .Q(state[8]) );
  DFFQX1TS \state_reg[6]  ( .D(nextstate[6]), .CK(clk), .Q(state[6]) );
  DFFQX1TS \state_reg[3]  ( .D(nextstate[3]), .CK(clk), .Q(state[3]) );
  CLKBUFX2TS U3 ( .A(sr_mp[0]), .Y(reg_ep) );
  CLKBUFX2TS U4 ( .A(sr_mq[0]), .Y(reg_eq) );
  OR3X2TS U5 ( .A(mux4[0]), .B(mux4[1]), .C(mux10), .Y(reg_ms) );
  AOI21X2TS U6 ( .A0(n499), .A1(n496), .B0(reset), .Y(reg_mc) );
  OAI211X2TS U7 ( .A0(reset), .A1(n596), .B0(n595), .C0(n594), .Y(mux14[1]) );
  CLKBUFX2TS U8 ( .A(reg_acc), .Y(mux1[0]) );
  NOR2X4TS U9 ( .A(reset), .B(n474), .Y(reg_r) );
  NOR2X4TS U10 ( .A(reset), .B(n546), .Y(reg_reg) );
  NOR2XLTS U11 ( .A(n525), .B(n146), .Y(n218) );
  NOR2XLTS U12 ( .A(n189), .B(n408), .Y(n232) );
  NOR2XLTS U13 ( .A(n503), .B(n408), .Y(n105) );
  NAND3XLTS U14 ( .A(state[1]), .B(state[3]), .C(n396), .Y(n14) );
  NAND3XLTS U15 ( .A(state[1]), .B(n514), .C(n401), .Y(n35) );
  AOI211XLTS U16 ( .A0(n572), .A1(n580), .B0(n218), .C0(n119), .Y(n465) );
  AOI211XLTS U17 ( .A0(n565), .A1(n582), .B0(n208), .C0(n2), .Y(n549) );
  NOR2XLTS U18 ( .A(n409), .B(n508), .Y(n13) );
  NOR2XLTS U19 ( .A(n484), .B(n82), .Y(n108) );
  NOR2XLTS U20 ( .A(n527), .B(n82), .Y(n107) );
  NAND3XLTS U21 ( .A(state[1]), .B(n401), .C(n515), .Y(n309) );
  NOR2XLTS U22 ( .A(n503), .B(n407), .Y(n449) );
  OAI211XLTS U23 ( .A0(n193), .A1(n367), .B0(n192), .C0(n191), .Y(n588) );
  OAI211XLTS U24 ( .A0(n407), .A1(n189), .B0(n211), .C0(n126), .Y(n313) );
  NOR2XLTS U25 ( .A(n293), .B(n82), .Y(n305) );
  NOR2XLTS U26 ( .A(n593), .B(n35), .Y(n172) );
  NOR2XLTS U27 ( .A(n527), .B(n367), .Y(n176) );
  NOR2XLTS U28 ( .A(n410), .B(n263), .Y(n473) );
  NOR2XLTS U29 ( .A(n513), .B(n138), .Y(n27) );
  NOR2XLTS U30 ( .A(n593), .B(n158), .Y(n28) );
  NOR2XLTS U31 ( .A(n407), .B(n367), .Y(n220) );
  AOI211XLTS U32 ( .A0(n577), .A1(n362), .B0(n227), .C0(n232), .Y(n370) );
  NOR2XLTS U33 ( .A(n101), .B(n407), .Y(n68) );
  OAI21XLTS U34 ( .A0(n260), .A1(n162), .B0(n580), .Y(n81) );
  NOR2XLTS U35 ( .A(n513), .B(n132), .Y(n227) );
  NAND3XLTS U36 ( .A(state[3]), .B(n396), .C(n590), .Y(n140) );
  NOR2XLTS U37 ( .A(n312), .B(n505), .Y(n279) );
  NOR2XLTS U38 ( .A(n525), .B(n585), .Y(n614) );
  CLKAND2X2TS U39 ( .A(n164), .B(n291), .Y(n208) );
  NOR2XLTS U40 ( .A(n312), .B(n157), .Y(n152) );
  NOR2XLTS U41 ( .A(n593), .B(n189), .Y(n103) );
  NOR2XLTS U42 ( .A(n10), .B(n446), .Y(n197) );
  NOR3BXLTS U43 ( .AN(n233), .B(n232), .C(n271), .Y(n236) );
  NOR2XLTS U44 ( .A(n312), .B(n82), .Y(n118) );
  NOR2XLTS U45 ( .A(n527), .B(n57), .Y(n119) );
  NOR2XLTS U46 ( .A(n304), .B(n289), .Y(n120) );
  OR2X1TS U47 ( .A(n391), .B(n9), .Y(n126) );
  NOR2XLTS U48 ( .A(n41), .B(n508), .Y(n125) );
  NOR2XLTS U49 ( .A(n590), .B(n288), .Y(n139) );
  NOR2XLTS U50 ( .A(n293), .B(n503), .Y(n109) );
  NOR2XLTS U51 ( .A(n12), .B(n304), .Y(n48) );
  OAI21XLTS U52 ( .A0(n557), .A1(n219), .B0(n15), .Y(n342) );
  AOI211XLTS U53 ( .A0(n203), .A1(n29), .B0(n176), .C0(n152), .Y(n257) );
  CLKAND2X2TS U54 ( .A(n610), .B(n611), .Y(n231) );
  NOR2XLTS U55 ( .A(n293), .B(n309), .Y(n356) );
  NOR2XLTS U56 ( .A(n304), .B(n146), .Y(n207) );
  NOR2XLTS U57 ( .A(n557), .B(n101), .Y(n460) );
  NAND3XLTS U58 ( .A(n291), .B(n577), .C(n415), .Y(n613) );
  NOR2XLTS U59 ( .A(n153), .B(n484), .Y(n314) );
  NOR2XLTS U60 ( .A(n409), .B(n513), .Y(n164) );
  NAND3XLTS U61 ( .A(state[6]), .B(state[7]), .C(state[5]), .Y(n45) );
  NAND3XLTS U62 ( .A(n465), .B(n549), .C(n464), .Y(n426) );
  NAND3XLTS U63 ( .A(state[6]), .B(state[5]), .C(n563), .Y(n7) );
  NOR2XLTS U64 ( .A(n397), .B(n416), .Y(n514) );
  OAI211XLTS U65 ( .A0(n309), .A1(n193), .B0(n23), .C0(n133), .Y(n604) );
  AOI211XLTS U66 ( .A0(n393), .A1(n362), .B0(n252), .C0(n251), .Y(n606) );
  NOR2XLTS U67 ( .A(n484), .B(n178), .Y(n93) );
  AOI211XLTS U68 ( .A0(n393), .A1(n32), .B0(n125), .C0(n108), .Y(n335) );
  NAND2BXLTS U69 ( .AN(n409), .B(n629), .Y(n263) );
  NAND3XLTS U70 ( .A(n577), .B(n415), .C(n531), .Y(n502) );
  NOR3XLTS U71 ( .A(n328), .B(n320), .C(n343), .Y(n457) );
  OAI21XLTS U72 ( .A0(n304), .A1(n263), .B0(n443), .Y(n454) );
  NAND4XLTS U73 ( .A(n299), .B(n335), .C(n128), .D(n34), .Y(n455) );
  AOI211XLTS U74 ( .A0(n33), .A1(n32), .B0(n107), .C0(n449), .Y(n34) );
  NOR2XLTS U75 ( .A(n7), .B(n397), .Y(n396) );
  INVX2TS U76 ( .A(state[8]), .Y(n397) );
  CLKAND2X2TS U77 ( .A(n302), .B(n301), .Y(n480) );
  AOI211XLTS U78 ( .A0(n580), .A1(n573), .B0(n194), .C0(n588), .Y(n478) );
  NOR2XLTS U79 ( .A(n189), .B(n312), .Y(n194) );
  NOR3XLTS U80 ( .A(n314), .B(n614), .C(n313), .Y(n475) );
  NOR2XLTS U81 ( .A(n312), .B(n439), .Y(n553) );
  OAI21XLTS U82 ( .A0(n294), .A1(n293), .B0(n438), .Y(n355) );
  NAND2BXLTS U83 ( .AN(n41), .B(n629), .Y(n620) );
  NAND4XLTS U84 ( .A(n352), .B(n192), .C(n257), .D(n248), .Y(n30) );
  NOR2XLTS U85 ( .A(n355), .B(n209), .Y(n98) );
  OAI21XLTS U86 ( .A0(n219), .A1(n484), .B0(n262), .Y(n226) );
  NOR2XLTS U87 ( .A(n152), .B(n162), .Y(n154) );
  NAND3XLTS U88 ( .A(n221), .B(n495), .C(n636), .Y(n166) );
  OAI21XLTS U89 ( .A0(n303), .A1(n525), .B0(n436), .Y(n209) );
  NAND3BXLTS U90 ( .AN(n241), .B(n357), .C(n624), .Y(n142) );
  AOI211XLTS U91 ( .A0(n435), .A1(n190), .B0(n109), .C0(n604), .Y(n24) );
  NAND4XLTS U92 ( .A(n257), .B(n606), .C(n256), .D(n255), .Y(n477) );
  NAND3XLTS U93 ( .A(n231), .B(n620), .C(n371), .Y(n328) );
  OAI211XLTS U94 ( .A0(n497), .A1(n555), .B0(n568), .C0(n613), .Y(n4) );
  INVX2TS U95 ( .A(state[2]), .Y(n569) );
  NOR2XLTS U96 ( .A(n7), .B(n10), .Y(n501) );
  NOR4BXLTS U97 ( .AN(n268), .B(n3), .C(n93), .D(n58), .Y(n568) );
  NOR2XLTS U98 ( .A(n469), .B(n138), .Y(n3) );
  INVX2TS U99 ( .A(state[1]), .Y(n590) );
  NOR2XLTS U100 ( .A(n455), .B(n454), .Y(n456) );
  INVX2TS U101 ( .A(state[0]), .Y(n422) );
  INVX2TS U102 ( .A(state[3]), .Y(n416) );
  INVX2TS U103 ( .A(state[5]), .Y(n559) );
  INVX2TS U104 ( .A(state[6]), .Y(n536) );
  NOR4BXLTS U105 ( .AN(n478), .B(n553), .C(n477), .D(n476), .Y(n479) );
  NAND4XLTS U106 ( .A(n475), .B(n550), .C(n474), .D(n599), .Y(n476) );
  NAND3XLTS U107 ( .A(n635), .B(n277), .C(n274), .Y(n184) );
  CLKBUFX2TS U108 ( .A(n56), .Y(reg_acc) );
  AO21X2TS U109 ( .A0(n471), .A1(n421), .B0(mux21[0]), .Y(reg_sum) );
  INVX2TS U110 ( .A(reset), .Y(n471) );
  NOR2XLTS U111 ( .A(state[1]), .B(state[8]), .Y(n417) );
  NAND2X1TS U112 ( .A(state[3]), .B(n417), .Y(n525) );
  NOR2XLTS U113 ( .A(state[6]), .B(state[7]), .Y(n489) );
  NAND2X1TS U114 ( .A(n489), .B(n559), .Y(n446) );
  NOR2X1TS U115 ( .A(n525), .B(n446), .Y(n630) );
  INVX2TS U116 ( .A(state[4]), .Y(n411) );
  NAND2X1TS U117 ( .A(state[2]), .B(state[0]), .Y(n526) );
  NOR2X1TS U118 ( .A(n411), .B(n526), .Y(n582) );
  NAND2X1TS U119 ( .A(n630), .B(n582), .Y(n546) );
  NAND2X1TS U120 ( .A(state[2]), .B(n422), .Y(n557) );
  NOR2X2TS U121 ( .A(state[4]), .B(n557), .Y(n577) );
  INVX2TS U122 ( .A(n577), .Y(n312) );
  NAND2X1TS U123 ( .A(state[3]), .B(n397), .Y(n584) );
  NOR2X1TS U124 ( .A(n590), .B(n584), .Y(n524) );
  INVX2TS U125 ( .A(n446), .Y(n401) );
  NAND2X1TS U126 ( .A(n524), .B(n401), .Y(n439) );
  INVX2TS U127 ( .A(n417), .Y(n264) );
  NOR2X1TS U128 ( .A(state[3]), .B(n264), .Y(n276) );
  NAND2X1TS U129 ( .A(n276), .B(n401), .Y(n101) );
  NOR2XLTS U130 ( .A(n397), .B(state[3]), .Y(n515) );
  NAND2X1TS U131 ( .A(n590), .B(n515), .Y(n9) );
  INVX2TS U132 ( .A(n9), .Y(n523) );
  NAND2X1TS U133 ( .A(n401), .B(n523), .Y(n367) );
  INVX2TS U134 ( .A(n367), .Y(n572) );
  NOR2X1TS U135 ( .A(state[2]), .B(state[4]), .Y(n631) );
  NAND2X1TS U136 ( .A(n631), .B(n422), .Y(n293) );
  INVX2TS U137 ( .A(n293), .Y(n580) );
  NOR3X1TS U138 ( .A(state[6]), .B(state[7]), .C(n559), .Y(n415) );
  NOR2X1TS U139 ( .A(state[2]), .B(n411), .Y(n253) );
  NAND2X1TS U140 ( .A(n253), .B(n422), .Y(n193) );
  INVX2TS U141 ( .A(n193), .Y(n203) );
  NAND2X1TS U142 ( .A(n415), .B(n203), .Y(n146) );
  NOR2X1TS U143 ( .A(n411), .B(n557), .Y(n190) );
  INVX2TS U144 ( .A(n190), .Y(n527) );
  INVX2TS U145 ( .A(n525), .Y(n291) );
  INVX2TS U146 ( .A(state[7]), .Y(n563) );
  NOR3X1TS U147 ( .A(state[6]), .B(state[5]), .C(n563), .Y(n111) );
  NAND2X1TS U148 ( .A(n291), .B(n111), .Y(n57) );
  INVX2TS U149 ( .A(n57), .Y(n565) );
  NAND2X1TS U150 ( .A(state[0]), .B(n415), .Y(n409) );
  INVX2TS U151 ( .A(n253), .Y(n513) );
  NOR2X1TS U152 ( .A(state[4]), .B(n569), .Y(n629) );
  INVX2TS U153 ( .A(n629), .Y(n504) );
  NOR2X1TS U154 ( .A(n7), .B(n9), .Y(n554) );
  NAND2X1TS U155 ( .A(state[0]), .B(n554), .Y(n132) );
  NAND2X1TS U156 ( .A(n631), .B(state[0]), .Y(n408) );
  OAI22X1TS U157 ( .A0(n504), .A1(n132), .B0(n367), .B1(n408), .Y(n2) );
  NAND2X1TS U158 ( .A(n554), .B(n577), .Y(n464) );
  INVX2TS U159 ( .A(n630), .Y(n497) );
  NAND2X1TS U160 ( .A(state[0]), .B(n569), .Y(n555) );
  NAND2X1TS U161 ( .A(n397), .B(n416), .Y(n556) );
  NOR2X1TS U162 ( .A(n590), .B(n556), .Y(n531) );
  NAND2X1TS U163 ( .A(state[2]), .B(state[4]), .Y(n508) );
  NAND2X1TS U164 ( .A(n531), .B(n13), .Y(n268) );
  INVX2TS U165 ( .A(n631), .Y(n469) );
  NAND2X1TS U166 ( .A(n396), .B(n416), .Y(n288) );
  NAND2X1TS U167 ( .A(state[0]), .B(n139), .Y(n138) );
  INVX2TS U168 ( .A(n582), .Y(n484) );
  INVX2TS U169 ( .A(n45), .Y(n482) );
  NAND2X1TS U170 ( .A(n524), .B(n482), .Y(n178) );
  INVX2TS U171 ( .A(n524), .Y(n304) );
  INVX2TS U172 ( .A(n111), .Y(n289) );
  NAND2X1TS U173 ( .A(state[0]), .B(n253), .Y(n407) );
  NOR2BX1TS U174 ( .AN(n120), .B(n407), .Y(n58) );
  NOR4X1TS U175 ( .A(n553), .B(n460), .C(n426), .D(n4), .Y(n659) );
  AOI22X1TS U176 ( .A0(n190), .A1(n120), .B0(n577), .B1(n139), .Y(n334) );
  INVX2TS U177 ( .A(n309), .Y(n435) );
  INVX2TS U178 ( .A(n408), .Y(n434) );
  AOI22X1TS U179 ( .A0(n577), .A1(n572), .B0(n435), .B1(n434), .Y(n635) );
  NOR3X1TS U180 ( .A(state[6]), .B(n563), .C(n559), .Y(n578) );
  NAND2X1TS U181 ( .A(n276), .B(n578), .Y(n249) );
  NAND2X1TS U182 ( .A(n249), .B(n140), .Y(n29) );
  INVX2TS U183 ( .A(n29), .Y(n294) );
  INVX2TS U184 ( .A(n138), .Y(n87) );
  AOI22X1TS U185 ( .A0(n629), .A1(n87), .B0(n120), .B1(n582), .Y(n438) );
  INVX2TS U186 ( .A(n415), .Y(n394) );
  NOR2X1TS U187 ( .A(n527), .B(n394), .Y(n290) );
  INVX2TS U188 ( .A(n290), .Y(n303) );
  NAND2X1TS U189 ( .A(n524), .B(n164), .Y(n436) );
  NAND2X1TS U190 ( .A(n635), .B(n98), .Y(n462) );
  NOR4BXLTS U191 ( .AN(n334), .B(n207), .C(n356), .D(n462), .Y(n658) );
  INVX2TS U192 ( .A(n276), .Y(n410) );
  NAND2X1TS U193 ( .A(n590), .B(n514), .Y(n10) );
  INVX2TS U194 ( .A(n197), .Y(n180) );
  INVX2TS U195 ( .A(n526), .Y(n402) );
  NAND2X1TS U196 ( .A(n402), .B(n411), .Y(n593) );
  INVX2TS U197 ( .A(n593), .Y(n626) );
  NAND2X1TS U198 ( .A(n626), .B(n435), .Y(n6) );
  OAI21XLTS U199 ( .A0(n203), .A1(n582), .B0(n572), .Y(n5) );
  OAI211XLTS U200 ( .A0(n407), .A1(n180), .B0(n6), .C0(n5), .Y(n175) );
  NAND2X1TS U201 ( .A(n578), .B(n291), .Y(n189) );
  NAND2X1TS U202 ( .A(n197), .B(n582), .Y(n211) );
  NAND2X1TS U203 ( .A(n111), .B(n434), .Y(n391) );
  NOR3XLTS U204 ( .A(n473), .B(n175), .C(n313), .Y(n70) );
  INVX2TS U205 ( .A(n14), .Y(n307) );
  NAND2X1TS U206 ( .A(state[0]), .B(n307), .Y(n41) );
  NAND2X1TS U207 ( .A(state[0]), .B(n501), .Y(n250) );
  INVX2TS U208 ( .A(n250), .Y(n254) );
  AOI22X1TS U209 ( .A0(state[4]), .A1(n254), .B0(n190), .B1(n554), .Y(n8) );
  OAI21XLTS U210 ( .A0(n469), .A1(n41), .B0(n8), .Y(n75) );
  NOR2XLTS U211 ( .A(n263), .B(n9), .Y(n205) );
  NOR2XLTS U212 ( .A(n10), .B(n391), .Y(n266) );
  NOR2XLTS U213 ( .A(n205), .B(n266), .Y(n155) );
  INVX2TS U214 ( .A(n407), .Y(n393) );
  NOR3X1TS U215 ( .A(state[7]), .B(state[5]), .C(n536), .Y(n579) );
  NAND2X1TS U216 ( .A(n276), .B(n579), .Y(n153) );
  INVX2TS U217 ( .A(n153), .Y(n165) );
  INVX2TS U218 ( .A(n13), .Y(n44) );
  NOR2XLTS U219 ( .A(n304), .B(n44), .Y(n311) );
  NAND2X1TS U220 ( .A(n579), .B(n291), .Y(n157) );
  AOI21X1TS U221 ( .A0(n293), .A1(n593), .B0(n157), .Y(n11) );
  AOI211XLTS U222 ( .A0(n393), .A1(n165), .B0(n311), .C0(n11), .Y(n65) );
  INVX2TS U223 ( .A(n101), .Y(n321) );
  NOR2XLTS U224 ( .A(n525), .B(n263), .Y(n77) );
  NOR2XLTS U225 ( .A(n593), .B(n439), .Y(n198) );
  AOI211XLTS U226 ( .A0(n402), .A1(n321), .B0(n77), .C0(n198), .Y(n340) );
  INVX2TS U227 ( .A(n439), .Y(n627) );
  INVX2TS U228 ( .A(n579), .Y(n12) );
  INVX2TS U229 ( .A(n48), .Y(n159) );
  NOR2XLTS U230 ( .A(n407), .B(n159), .Y(n366) );
  INVX2TS U231 ( .A(n531), .Y(n483) );
  NOR2XLTS U232 ( .A(n263), .B(n483), .Y(n642) );
  AOI211XLTS U233 ( .A0(n582), .A1(n627), .B0(n366), .C0(n642), .Y(n270) );
  NAND4XLTS U234 ( .A(n155), .B(n65), .C(n340), .D(n270), .Y(n22) );
  OAI22X1TS U235 ( .A0(n411), .A1(n249), .B0(n189), .B1(n312), .Y(n84) );
  AOI22X1TS U236 ( .A0(n291), .A1(n13), .B0(n524), .B1(n290), .Y(n64) );
  AOI22X1TS U237 ( .A0(n626), .A1(n572), .B0(n577), .B1(n435), .Y(n173) );
  NAND2X1TS U238 ( .A(n153), .B(n180), .Y(n362) );
  AOI22X1TS U239 ( .A0(n580), .A1(n362), .B0(n577), .B1(n29), .Y(n302) );
  NAND2X1TS U240 ( .A(n578), .B(n531), .Y(n82) );
  OAI22X1TS U241 ( .A0(n469), .A1(n250), .B0(n293), .B1(n14), .Y(n76) );
  NOR2X1TS U242 ( .A(n446), .B(n483), .Y(n625) );
  INVX2TS U243 ( .A(n625), .Y(n219) );
  NAND2X1TS U244 ( .A(n524), .B(n415), .Y(n505) );
  AOI21X1TS U245 ( .A0(n203), .A1(n321), .B0(n279), .Y(n15) );
  OAI22X1TS U246 ( .A0(n439), .A1(n555), .B0(n249), .B1(n408), .Y(n16) );
  NOR4XLTS U247 ( .A(n305), .B(n76), .C(n342), .D(n16), .Y(n17) );
  AND4X1TS U248 ( .A(n64), .B(n173), .C(n302), .D(n17), .Y(n458) );
  NAND4XLTS U249 ( .A(state[6]), .B(state[7]), .C(n276), .D(n434), .Y(n18) );
  NOR2XLTS U250 ( .A(state[5]), .B(n18), .Y(n364) );
  NOR2XLTS U251 ( .A(n484), .B(n157), .Y(n271) );
  NOR2XLTS U252 ( .A(n364), .B(n271), .Y(n326) );
  NOR3XLTS U253 ( .A(state[2]), .B(state[0]), .C(n439), .Y(n361) );
  NOR2XLTS U254 ( .A(n469), .B(n409), .Y(n163) );
  NAND2X1TS U255 ( .A(n524), .B(n163), .Y(n494) );
  INVX2TS U256 ( .A(n494), .Y(n643) );
  AOI22X1TS U257 ( .A0(n203), .A1(n120), .B0(n531), .B1(n290), .Y(n19) );
  NAND2X1TS U258 ( .A(n580), .B(n139), .Y(n357) );
  OAI211XLTS U259 ( .A0(n178), .A1(n527), .B0(n19), .C0(n357), .Y(n331) );
  NAND2X1TS U260 ( .A(n276), .B(n163), .Y(n552) );
  NAND2BXLTS U261 ( .AN(n331), .B(n552), .Y(n430) );
  NOR4XLTS U262 ( .A(n321), .B(n361), .C(n643), .D(n430), .Y(n20) );
  NAND4BXLTS U263 ( .AN(n84), .B(n458), .C(n326), .D(n20), .Y(n21) );
  NOR4BXLTS U264 ( .AN(n70), .B(n75), .C(n22), .D(n21), .Y(n657) );
  OAI22X1TS U265 ( .A0(n508), .A1(n132), .B0(n408), .B1(n157), .Y(n31) );
  NAND2X1TS U266 ( .A(state[1]), .B(n396), .Y(n25) );
  NAND2X1TS U267 ( .A(n578), .B(n524), .Y(n503) );
  INVX2TS U268 ( .A(n503), .Y(n85) );
  AOI22X1TS U269 ( .A0(n580), .A1(n48), .B0(n577), .B1(n85), .Y(n23) );
  NAND2X1TS U270 ( .A(n190), .B(n139), .Y(n133) );
  AOI32X1TS U271 ( .A0(n25), .A1(n24), .A2(n82), .B0(n193), .B1(n24), .Y(n26)
         );
  NAND2X1TS U272 ( .A(n579), .B(n531), .Y(n158) );
  NAND2X1TS U273 ( .A(n35), .B(n158), .Y(n32) );
  OAI32X1TS U274 ( .A0(n26), .A1(n48), .A2(n32), .B0(n577), .B1(n26), .Y(n352)
         );
  NOR4XLTS U275 ( .A(n28), .B(n105), .C(n172), .D(n27), .Y(n192) );
  AOI22X1TS U276 ( .A0(n190), .A1(n29), .B0(n203), .B1(n362), .Y(n248) );
  NOR4XLTS U277 ( .A(n103), .B(n220), .C(n31), .D(n30), .Y(n299) );
  NOR4XLTS U278 ( .A(state[3]), .B(n397), .C(n590), .D(n391), .Y(n448) );
  AOI21X1TS U279 ( .A0(n190), .A1(n307), .B0(n448), .Y(n128) );
  NAND2X1TS U280 ( .A(n193), .B(n484), .Y(n33) );
  INVX2TS U281 ( .A(n158), .Y(n162) );
  NAND2X1TS U282 ( .A(n162), .B(n434), .Y(n610) );
  INVX2TS U283 ( .A(n82), .Y(n500) );
  NAND2X1TS U284 ( .A(n626), .B(n500), .Y(n611) );
  INVX2TS U285 ( .A(n35), .Y(n260) );
  NAND2X1TS U286 ( .A(n260), .B(n434), .Y(n371) );
  OAI22X1TS U287 ( .A0(n557), .A1(n497), .B0(n410), .B1(n146), .Y(n320) );
  INVX2TS U288 ( .A(n189), .Y(n112) );
  AOI22X1TS U289 ( .A0(n580), .A1(n112), .B0(n165), .B1(n626), .Y(n196) );
  AOI22X1TS U290 ( .A0(n554), .A1(n203), .B0(n626), .B1(n197), .Y(n649) );
  NOR2BX1TS U291 ( .AN(n81), .B(n118), .Y(n244) );
  AND4X1TS U292 ( .A(n196), .B(n649), .C(n370), .D(n244), .Y(n36) );
  NAND2X1TS U293 ( .A(n307), .B(n577), .Y(n277) );
  NAND2X1TS U294 ( .A(n36), .B(n277), .Y(n343) );
  NAND2X1TS U295 ( .A(n203), .B(n625), .Y(n597) );
  NOR2X1TS U296 ( .A(n293), .B(n394), .Y(n275) );
  NAND2X1TS U297 ( .A(n524), .B(n275), .Y(n598) );
  AND3X1TS U298 ( .A(n546), .B(n597), .C(n598), .Y(n318) );
  NOR2XLTS U299 ( .A(n593), .B(n497), .Y(n461) );
  INVX2TS U300 ( .A(n555), .Y(n530) );
  NAND2X1TS U301 ( .A(n625), .B(n530), .Y(n599) );
  INVX2TS U302 ( .A(n599), .Y(n459) );
  NOR2XLTS U303 ( .A(n461), .B(n459), .Y(n596) );
  NAND2X1TS U304 ( .A(n276), .B(n415), .Y(n592) );
  NOR2XLTS U305 ( .A(n407), .B(n592), .Y(n67) );
  INVX2TS U306 ( .A(n67), .Y(n539) );
  NAND4XLTS U307 ( .A(n457), .B(n318), .C(n596), .D(n539), .Y(n452) );
  INVX2TS U308 ( .A(n157), .Y(n573) );
  AOI22X1TS U309 ( .A0(n580), .A1(n554), .B0(n203), .B1(n565), .Y(n38) );
  NOR2XLTS U310 ( .A(n525), .B(n45), .Y(n37) );
  NAND2X1TS U311 ( .A(n190), .B(n37), .Y(n150) );
  NAND2X1TS U312 ( .A(n276), .B(n290), .Y(n272) );
  NAND3XLTS U313 ( .A(n38), .B(n150), .C(n272), .Y(n330) );
  AOI211XLTS U314 ( .A0(n393), .A1(n573), .B0(n314), .C0(n330), .Y(n39) );
  NAND2X1TS U315 ( .A(n580), .B(n625), .Y(n322) );
  NAND4XLTS U316 ( .A(n39), .B(n471), .C(n82), .D(n322), .Y(n55) );
  OAI22X1TS U317 ( .A0(n250), .A1(n504), .B0(n593), .B1(n249), .Y(n40) );
  AOI21X1TS U318 ( .A0(n434), .A1(n362), .B0(n40), .Y(n301) );
  NOR2XLTS U319 ( .A(n41), .B(n513), .Y(n96) );
  NOR2XLTS U320 ( .A(n508), .B(n138), .Y(n95) );
  NOR2XLTS U321 ( .A(n408), .B(n159), .Y(n60) );
  AOI21X1TS U322 ( .A0(n85), .A1(n626), .B0(n60), .Y(n238) );
  NAND2X1TS U323 ( .A(n393), .B(n435), .Y(n42) );
  NAND4BXLTS U324 ( .AN(n95), .B(n238), .C(n502), .D(n42), .Y(n603) );
  AOI22X1TS U325 ( .A0(n630), .A1(n203), .B0(n531), .B1(n164), .Y(n43) );
  NAND2X1TS U326 ( .A(n531), .B(n275), .Y(n474) );
  OAI211XLTS U327 ( .A0(n309), .A1(n484), .B0(n43), .C0(n474), .Y(n230) );
  INVX2TS U328 ( .A(n514), .Y(n528) );
  NOR3XLTS U329 ( .A(n528), .B(n527), .C(n446), .Y(n183) );
  NAND3XLTS U330 ( .A(n580), .B(n111), .C(n515), .Y(n123) );
  INVX2TS U331 ( .A(n584), .Y(n560) );
  NAND3XLTS U332 ( .A(n578), .B(n560), .C(n203), .Y(n121) );
  INVX2TS U333 ( .A(n556), .Y(n507) );
  NAND2X1TS U334 ( .A(n579), .B(n507), .Y(n445) );
  OR2X1TS U335 ( .A(n445), .B(n527), .Y(n145) );
  NAND4BXLTS U336 ( .AN(n183), .B(n123), .C(n121), .D(n145), .Y(n545) );
  AOI21X1TS U337 ( .A0(n291), .A1(n163), .B0(n545), .Y(n297) );
  NOR2XLTS U338 ( .A(n410), .B(n44), .Y(n267) );
  NOR3XLTS U339 ( .A(n525), .B(n484), .C(n45), .Y(n59) );
  INVX2TS U340 ( .A(n59), .Y(n212) );
  NOR2XLTS U341 ( .A(n469), .B(n132), .Y(n66) );
  INVX2TS U342 ( .A(n66), .Y(n46) );
  OAI211XLTS U343 ( .A0(n57), .A1(n407), .B0(n212), .C0(n46), .Y(n412) );
  NOR2XLTS U344 ( .A(n267), .B(n412), .Y(n52) );
  NOR2XLTS U345 ( .A(n593), .B(n159), .Y(n61) );
  NOR2XLTS U346 ( .A(n527), .B(n439), .Y(n182) );
  AOI211XLTS U347 ( .A0(n275), .A1(n417), .B0(n61), .C0(n182), .Y(n51) );
  NOR2XLTS U348 ( .A(n483), .B(n146), .Y(n124) );
  INVX2TS U349 ( .A(n592), .Y(n317) );
  AO22XLTS U350 ( .A0(n577), .A1(n317), .B0(n531), .B1(n163), .Y(n300) );
  AOI22X1TS U351 ( .A0(n190), .A1(n112), .B0(n523), .B1(n275), .Y(n47) );
  NAND3XLTS U352 ( .A(n577), .B(n111), .C(n523), .Y(n122) );
  OAI211XLTS U353 ( .A0(n157), .A1(n193), .B0(n47), .C0(n122), .Y(n544) );
  NAND2X1TS U354 ( .A(n500), .B(n393), .Y(n233) );
  NAND2X1TS U355 ( .A(n203), .B(n48), .Y(n149) );
  OAI211XLTS U356 ( .A0(n497), .A1(n293), .B0(n233), .C0(n149), .Y(n49) );
  NOR4XLTS U357 ( .A(n124), .B(n300), .C(n544), .D(n49), .Y(n50) );
  NAND4XLTS U358 ( .A(n297), .B(n52), .C(n51), .D(n50), .Y(n53) );
  NOR4XLTS U359 ( .A(n96), .B(n603), .C(n230), .D(n53), .Y(n347) );
  AOI21X1TS U360 ( .A0(n625), .A1(n402), .B0(n68), .Y(n443) );
  AOI21X1TS U361 ( .A0(n321), .A1(n434), .B0(n454), .Y(n298) );
  NAND3XLTS U362 ( .A(n301), .B(n347), .C(n298), .Y(n54) );
  NOR4XLTS U363 ( .A(n455), .B(n452), .C(n55), .D(n54), .Y(n656) );
  NAND4XLTS U364 ( .A(n659), .B(n658), .C(n657), .D(n656), .Y(n660) );
  NOR3XLTS U365 ( .A(reset), .B(n407), .C(n157), .Y(n56) );
  NAND2X1TS U366 ( .A(N2139), .B(ms0_24), .Y(n383) );
  OAI21XLTS U367 ( .A0(N2139), .A1(ms0_24), .B0(n383), .Y(n644) );
  AOI32X1TS U368 ( .A0(n497), .A1(n268), .A2(n57), .B0(n407), .B1(n268), .Y(
        n224) );
  AOI211XLTS U369 ( .A0(n434), .A1(n630), .B0(n58), .C0(n224), .Y(n74) );
  AOI31XLTS U370 ( .A0(state[1]), .A1(n275), .A2(n397), .B0(n59), .Y(n63) );
  INVX2TS U371 ( .A(mq47), .Y(n360) );
  AOI211XLTS U372 ( .A0(n207), .A1(n360), .B0(n61), .C0(n60), .Y(n62) );
  NAND4XLTS U373 ( .A(n65), .B(n64), .C(n63), .D(n62), .Y(n168) );
  INVX2TS U374 ( .A(mode[2]), .Y(n641) );
  NAND2X1TS U375 ( .A(mode[0]), .B(n641), .Y(n359) );
  INVX2TS U376 ( .A(mode[0]), .Y(n639) );
  NAND2X1TS U377 ( .A(mode[2]), .B(n639), .Y(n195) );
  AOI21X1TS U378 ( .A0(n359), .A1(n195), .B0(mode[1]), .Y(n71) );
  NOR4BXLTS U379 ( .AN(n552), .B(n68), .C(n67), .D(n66), .Y(n69) );
  OAI211XLTS U380 ( .A0(n71), .A1(n322), .B0(n70), .C0(n69), .Y(n72) );
  AOI211XLTS U381 ( .A0(sumor), .A1(n330), .B0(n168), .C0(n72), .Y(n73) );
  NAND4XLTS U382 ( .A(n173), .B(n74), .C(n73), .D(n277), .Y(n100) );
  NOR2XLTS U383 ( .A(n76), .B(n75), .Y(n136) );
  NOR4XLTS U384 ( .A(n279), .B(n461), .C(n553), .D(n77), .Y(n78) );
  OAI211XLTS U385 ( .A0(n196), .A1(N2152), .B0(n136), .C0(n78), .Y(n623) );
  OAI22X1TS U386 ( .A0(N2152), .A1(n649), .B0(n334), .B1(mq47), .Y(n91) );
  OAI22X1TS U387 ( .A0(n527), .A1(n219), .B0(n484), .B1(n101), .Y(n79) );
  NOR2XLTS U388 ( .A(n267), .B(n79), .Y(n202) );
  AOI22X1TS U389 ( .A0(n626), .A1(n321), .B0(n577), .B1(n625), .Y(n80) );
  NAND4XLTS U390 ( .A(n81), .B(n202), .C(n80), .D(n464), .Y(n90) );
  AOI21X1TS U391 ( .A0(n469), .A1(n407), .B0(n82), .Y(n83) );
  AOI211XLTS U392 ( .A0(n626), .A1(n85), .B0(n84), .C0(n83), .Y(n106) );
  OAI22X1TS U393 ( .A0(ms0_23), .A1(n502), .B0(n249), .B1(n408), .Y(n86) );
  AOI211XLTS U394 ( .A0(n87), .A1(n631), .B0(n314), .C0(n86), .Y(n88) );
  OAI211XLTS U395 ( .A0(n635), .A1(N2131), .B0(n106), .C0(n88), .Y(n89) );
  NOR4XLTS U396 ( .A(n623), .B(n91), .C(n90), .D(n89), .Y(n382) );
  AOI22X1TS U397 ( .A0(mq47), .A1(n361), .B0(n366), .B1(r31), .Y(n92) );
  OAI211XLTS U398 ( .A0(n155), .A1(comp2_g), .B0(n465), .C0(n92), .Y(n336) );
  AOI21X1TS U399 ( .A0(n435), .A1(state[4]), .B0(n93), .Y(n187) );
  AOI21X1TS U400 ( .A0(n356), .A1(n360), .B0(n118), .Y(n637) );
  OAI211XLTS U401 ( .A0(N2152), .A1(n370), .B0(n187), .C0(n637), .Y(n94) );
  NOR4XLTS U402 ( .A(n96), .B(n95), .C(n336), .D(n94), .Y(n97) );
  OAI211XLTS U403 ( .A0(N2131), .A1(n98), .B0(n382), .C0(n97), .Y(n99) );
  AOI211XLTS U404 ( .A0(n328), .A1(n644), .B0(n100), .C0(n99), .Y(n102) );
  NOR3X1TS U405 ( .A(reset), .B(n101), .C(n408), .Y(mux21[0]) );
  NOR2XLTS U406 ( .A(reg_reg), .B(mux21[0]), .Y(n602) );
  AOI31XLTS U407 ( .A0(n102), .A1(n299), .A2(n602), .B0(reset), .Y(N2446) );
  NOR2XLTS U408 ( .A(n312), .B(n503), .Y(n104) );
  AOI211XLTS U409 ( .A0(n500), .A1(n203), .B0(n104), .C0(n103), .Y(n201) );
  NAND2BXLTS U410 ( .AN(n105), .B(n201), .Y(n372) );
  NAND4XLTS U411 ( .A(n106), .B(n212), .C(n611), .D(n150), .Y(n117) );
  NOR2XLTS U412 ( .A(n189), .B(n407), .Y(n110) );
  NOR4XLTS U413 ( .A(n110), .B(n109), .C(n108), .D(n107), .Y(n222) );
  NOR2XLTS U414 ( .A(n584), .B(n484), .Y(n481) );
  AOI22X1TS U415 ( .A0(n111), .A1(n481), .B0(n205), .B1(comp2_g), .Y(n115) );
  INVX2TS U416 ( .A(n249), .Y(n628) );
  AOI211XLTS U417 ( .A0(n112), .A1(n631), .B0(n628), .C0(n449), .Y(n114) );
  NAND2X1TS U418 ( .A(n190), .B(n120), .Y(n113) );
  NAND4XLTS U419 ( .A(n222), .B(n115), .C(n114), .D(n113), .Y(n116) );
  NOR4XLTS U420 ( .A(n118), .B(n372), .C(n117), .D(n116), .Y(n281) );
  AO21XLTS U421 ( .A0(n120), .A1(n253), .B0(n119), .Y(n204) );
  AOI32X1TS U422 ( .A0(n189), .A1(n121), .A2(n497), .B0(n527), .B1(n121), .Y(
        n167) );
  AOI211XLTS U423 ( .A0(n253), .A1(n565), .B0(n204), .C0(n167), .Y(n131) );
  NAND3BXLTS U424 ( .AN(n124), .B(n123), .C(n122), .Y(n171) );
  AOI21X1TS U425 ( .A0(n139), .A1(n203), .B0(n125), .Y(n127) );
  NAND3XLTS U426 ( .A(n128), .B(n127), .C(n126), .Y(n186) );
  OAI2BB2XLTS U427 ( .B0(N2139), .B1(n277), .A0N(comp2_g), .A1N(n364), .Y(n129) );
  NOR3XLTS U428 ( .A(n171), .B(n186), .C(n129), .Y(n130) );
  AOI31XLTS U429 ( .A0(n281), .A1(n131), .A2(n130), .B0(reset), .Y(N2452) );
  NAND2X1TS U430 ( .A(n138), .B(n132), .Y(n144) );
  INVX2TS U431 ( .A(n508), .Y(n571) );
  AOI22X1TS U432 ( .A0(n307), .A1(n253), .B0(n571), .B1(n144), .Y(n134) );
  NAND2X1TS U433 ( .A(n134), .B(n133), .Y(n215) );
  INVX2TS U434 ( .A(n554), .Y(n135) );
  NAND2X1TS U435 ( .A(n136), .B(n135), .Y(n143) );
  NAND2X1TS U436 ( .A(n254), .B(n629), .Y(n137) );
  OAI211XLTS U437 ( .A0(n140), .A1(n312), .B0(n620), .C0(n137), .Y(n241) );
  OAI22X1TS U438 ( .A0(n411), .A1(n140), .B0(n513), .B1(n138), .Y(n354) );
  OAI2BB2XLTS U439 ( .B0(n293), .B1(n140), .A0N(n577), .A1N(n139), .Y(n141) );
  AOI211XLTS U440 ( .A0(n629), .A1(n144), .B0(n354), .C0(n141), .Y(n624) );
  NOR4XLTS U441 ( .A(n144), .B(n215), .C(n143), .D(n142), .Y(n282) );
  OA21XLTS U442 ( .A0(n157), .A1(n193), .B0(n145), .Y(n540) );
  NOR2XLTS U443 ( .A(n410), .B(n146), .Y(n148) );
  INVX2TS U444 ( .A(n597), .Y(n147) );
  AOI211XLTS U445 ( .A0(n630), .A1(n577), .B0(n148), .C0(n147), .Y(n151) );
  NAND4XLTS U446 ( .A(n540), .B(n151), .C(n150), .D(n149), .Y(n214) );
  INVX2TS U447 ( .A(comp2_g), .Y(n363) );
  OAI211XLTS U448 ( .A0(n155), .A1(n363), .B0(n154), .C0(n153), .Y(n156) );
  AOI211XLTS U449 ( .A0(N2131), .A1(n209), .B0(n214), .C0(n156), .Y(n170) );
  NOR2XLTS U450 ( .A(n408), .B(n157), .Y(n161) );
  AOI21X1TS U451 ( .A0(n312), .A1(n513), .B0(n158), .Y(n369) );
  INVX2TS U452 ( .A(N2139), .Y(n344) );
  OAI22X1TS U453 ( .A0(n159), .A1(state[4]), .B0(n344), .B1(n277), .Y(n160) );
  NOR4XLTS U454 ( .A(n314), .B(n161), .C(n369), .D(n160), .Y(n243) );
  AOI22X1TS U455 ( .A0(n291), .A1(n163), .B0(n162), .B1(n582), .Y(n221) );
  NAND2X1TS U456 ( .A(n531), .B(n164), .Y(n495) );
  AOI22X1TS U457 ( .A0(n165), .A1(n577), .B0(n271), .B1(n363), .Y(n636) );
  NOR4BXLTS U458 ( .AN(n243), .B(n168), .C(n167), .D(n166), .Y(n169) );
  AOI31XLTS U459 ( .A0(n282), .A1(n170), .A2(n169), .B0(reset), .Y(N2451) );
  AOI211XLTS U460 ( .A0(n260), .A1(n580), .B0(n172), .C0(n171), .Y(n177) );
  AOI32X1TS U461 ( .A0(n469), .A1(n173), .A2(n193), .B0(n180), .B1(n173), .Y(
        n174) );
  NOR4BXLTS U462 ( .AN(n177), .B(n176), .C(n175), .D(n174), .Y(n618) );
  NOR2XLTS U463 ( .A(n527), .B(n178), .Y(n179) );
  AOI211XLTS U464 ( .A0(n266), .A1(comp2_g), .B0(n260), .C0(n179), .Y(n181) );
  INVX2TS U465 ( .A(n356), .Y(n333) );
  NAND4XLTS U466 ( .A(n181), .B(n180), .C(n367), .D(n333), .Y(n185) );
  AOI211XLTS U467 ( .A0(n275), .A1(n523), .B0(n183), .C0(n182), .Y(n274) );
  NOR4BXLTS U468 ( .AN(n187), .B(n186), .C(n185), .D(n184), .Y(n188) );
  AOI31XLTS U469 ( .A0(n282), .A1(n618), .A2(n188), .B0(reset), .Y(N2453) );
  NAND2X1TS U470 ( .A(n190), .B(n554), .Y(n191) );
  NOR2XLTS U471 ( .A(reset), .B(n478), .Y(ssr_ms0[1]) );
  INVX2TS U472 ( .A(N2152), .Y(n648) );
  OR2X1TS U473 ( .A(mode[1]), .B(n322), .Y(n638) );
  OAI22X1TS U474 ( .A0(n196), .A1(n648), .B0(n638), .B1(n195), .Y(n247) );
  AOI22X1TS U475 ( .A0(n577), .A1(n197), .B0(n625), .B1(n393), .Y(n200) );
  AOI21X1TS U476 ( .A0(n321), .A1(state[4]), .B0(n198), .Y(n199) );
  NAND4XLTS U477 ( .A(n202), .B(n201), .C(n200), .D(n199), .Y(n246) );
  OAI32X1TS U478 ( .A0(n364), .A1(n627), .A2(n565), .B0(n203), .B1(n364), .Y(
        n229) );
  NAND2X1TS U479 ( .A(n312), .B(n513), .Y(n206) );
  AOI211XLTS U480 ( .A0(n260), .A1(n206), .B0(n205), .C0(n204), .Y(n217) );
  INVX2TS U481 ( .A(n207), .Y(n332) );
  INVX2TS U482 ( .A(N2131), .Y(n634) );
  AOI21X1TS U483 ( .A0(n634), .A1(n209), .B0(n208), .Y(n210) );
  OAI21XLTS U484 ( .A0(n360), .A1(n332), .B0(n210), .Y(n286) );
  NAND4BXLTS U485 ( .AN(n449), .B(n212), .C(n211), .D(n546), .Y(n213) );
  NOR4XLTS U486 ( .A(n215), .B(n286), .C(n214), .D(n213), .Y(n216) );
  OAI211XLTS U487 ( .A0(n439), .A1(n407), .B0(n217), .C0(n216), .Y(n381) );
  AOI21X1TS U488 ( .A0(n290), .A1(n531), .B0(n218), .Y(n262) );
  AOI21X1TS U489 ( .A0(n435), .A1(state[4]), .B0(n220), .Y(n223) );
  NAND4BXLTS U490 ( .AN(n224), .B(n223), .C(n222), .D(n221), .Y(n225) );
  NOR4XLTS U491 ( .A(n227), .B(n381), .C(n226), .D(n225), .Y(n228) );
  NAND4BXLTS U492 ( .AN(n230), .B(n229), .C(n228), .D(n598), .Y(n653) );
  NOR2XLTS U493 ( .A(N2139), .B(ms0_24), .Y(n612) );
  INVX2TS U494 ( .A(n612), .Y(n619) );
  INVX2TS U495 ( .A(n322), .Y(n259) );
  NAND2X1TS U496 ( .A(n259), .B(mode[1]), .Y(n640) );
  OAI22X1TS U497 ( .A0(n231), .A1(n619), .B0(n640), .B1(n359), .Y(n240) );
  INVX2TS U498 ( .A(n371), .Y(n645) );
  NOR2XLTS U499 ( .A(n304), .B(n263), .Y(n265) );
  AOI21X1TS U500 ( .A0(n645), .A1(n383), .B0(n265), .Y(n237) );
  INVX2TS U501 ( .A(n272), .Y(n234) );
  AOI21X1TS U502 ( .A0(n363), .A1(n266), .B0(n234), .Y(n235) );
  NAND4XLTS U503 ( .A(n238), .B(n237), .C(n236), .D(n235), .Y(n239) );
  NOR4XLTS U504 ( .A(n653), .B(n241), .C(n240), .D(n239), .Y(n242) );
  OAI211XLTS U505 ( .A0(N2139), .A1(n244), .B0(n243), .C0(n242), .Y(n245) );
  NOR4BXLTS U506 ( .AN(n649), .B(n247), .C(n246), .D(n245), .Y(n258) );
  INVX2TS U507 ( .A(n248), .Y(n252) );
  OAI22X1TS U508 ( .A0(n250), .A1(n508), .B0(n484), .B1(n249), .Y(n251) );
  AOI22X1TS U509 ( .A0(n582), .A1(n572), .B0(n393), .B1(n628), .Y(n256) );
  AOI22X1TS U510 ( .A0(n254), .A1(n253), .B0(n626), .B1(n573), .Y(n255) );
  NAND2X1TS U511 ( .A(n477), .B(n471), .Y(n608) );
  INVX2TS U512 ( .A(n608), .Y(mux20[0]) );
  NOR2XLTS U513 ( .A(mux20[0]), .B(ssr_ms0[1]), .Y(n316) );
  NOR2X1TS U514 ( .A(reset), .B(n539), .Y(mux21[1]) );
  INVX2TS U515 ( .A(mux21[1]), .Y(n595) );
  OAI211XLTS U516 ( .A0(reset), .A1(n258), .B0(n316), .C0(n595), .Y(N2449) );
  AOI22X1TS U517 ( .A0(n260), .A1(n582), .B0(n259), .B1(mode[2]), .Y(n261) );
  OAI211XLTS U518 ( .A0(n264), .A1(n263), .B0(n262), .C0(n261), .Y(n285) );
  NOR4BXLTS U519 ( .AN(n268), .B(n267), .C(n266), .D(n265), .Y(n269) );
  OAI211XLTS U520 ( .A0(mode[0]), .A1(n640), .B0(n270), .C0(n269), .Y(n284) );
  INVX2TS U521 ( .A(n275), .Y(n585) );
  AOI211XLTS U522 ( .A0(n271), .A1(comp2_g), .B0(n643), .C0(n300), .Y(n273) );
  NAND4XLTS U523 ( .A(n274), .B(n273), .C(n272), .D(n613), .Y(n353) );
  NAND2X1TS U524 ( .A(n276), .B(n275), .Y(n442) );
  OAI211XLTS U525 ( .A0(n344), .A1(n277), .B0(n502), .C0(n442), .Y(n278) );
  NOR4XLTS U526 ( .A(n279), .B(n614), .C(n353), .D(n278), .Y(n280) );
  NAND3XLTS U527 ( .A(n282), .B(n281), .C(n280), .Y(n283) );
  NOR4XLTS U528 ( .A(n286), .B(n285), .C(n284), .D(n283), .Y(n287) );
  AOI31XLTS U529 ( .A0(n287), .A1(n552), .A2(n539), .B0(reset), .Y(N2450) );
  OAI32X1TS U530 ( .A0(n411), .A1(n584), .A2(n289), .B0(state[4]), .B1(n288), 
        .Y(n490) );
  AOI33XLTS U531 ( .A0(n559), .A1(n411), .A2(n515), .B0(state[5]), .B1(n560), 
        .B2(state[4]), .Y(n486) );
  INVX2TS U532 ( .A(n486), .Y(n535) );
  NAND3XLTS U533 ( .A(n569), .B(n536), .C(n535), .Y(n561) );
  AOI2BB2XLTS U534 ( .B0(state[2]), .B1(n490), .A0N(state[7]), .A1N(n561), .Y(
        n387) );
  AOI22X1TS U535 ( .A0(n291), .A1(n290), .B0(n577), .B1(n572), .Y(n292) );
  OAI32X1TS U536 ( .A0(reset), .A1(n294), .A2(n293), .B0(n292), .B1(reset), 
        .Y(mux7) );
  INVX2TS U537 ( .A(mux7), .Y(n432) );
  OAI31X1TS U538 ( .A0(reset), .A1(n387), .A2(n590), .B0(n432), .Y(reg_sp) );
  AOI21X1TS U539 ( .A0(n659), .A1(n458), .B0(reset), .Y(sr_mq[0]) );
  AOI21X1TS U540 ( .A0(n299), .A1(n658), .B0(reset), .Y(sr_mp[0]) );
  NOR2X1TS U541 ( .A(reset), .B(n297), .Y(mux2[0]) );
  OAI31X1TS U542 ( .A0(reset), .A1(n469), .A2(n505), .B0(n595), .Y(mux22) );
  INVX2TS U543 ( .A(mux22), .Y(n601) );
  OAI31X1TS U544 ( .A0(reset), .A1(n526), .A2(n497), .B0(n601), .Y(mux13[0])
         );
  AO21XLTS U545 ( .A0(n471), .A1(n459), .B0(mux13[0]), .Y(mux3[1]) );
  NOR2XLTS U546 ( .A(reset), .B(n298), .Y(rf_wa[1]) );
  AOI21X1TS U547 ( .A0(n659), .A1(n658), .B0(reset), .Y(mux17[2]) );
  NOR2XLTS U548 ( .A(reset), .B(n299), .Y(sr_mp[1]) );
  NOR2XLTS U549 ( .A(reset), .B(n458), .Y(sr_mq[1]) );
  NAND2X1TS U550 ( .A(n471), .B(n300), .Y(n431) );
  INVX2TS U551 ( .A(n431), .Y(counterii[1]) );
  NOR2XLTS U552 ( .A(n304), .B(n303), .Y(n306) );
  AOI211XLTS U553 ( .A0(n307), .A1(n631), .B0(n306), .C0(n305), .Y(n308) );
  OAI31X1TS U554 ( .A0(state[4]), .A1(n569), .A2(n309), .B0(n308), .Y(n310) );
  AOI211XLTS U555 ( .A0(n434), .A1(n500), .B0(n311), .C0(n310), .Y(n346) );
  NAND2X1TS U556 ( .A(n480), .B(n346), .Y(n466) );
  NOR3XLTS U557 ( .A(reset), .B(n312), .C(n592), .Y(mux4[0]) );
  NOR2XLTS U558 ( .A(reset), .B(n475), .Y(mux12[0]) );
  AOI211XLTS U559 ( .A0(n471), .A1(n466), .B0(mux4[0]), .C0(mux12[0]), .Y(n315) );
  NAND2X1TS U560 ( .A(n316), .B(n315), .Y(ssr_ms0[0]) );
  NOR2XLTS U561 ( .A(reset), .B(n495), .Y(n319) );
  AOI211XLTS U562 ( .A0(n582), .A1(n317), .B0(n331), .C0(n412), .Y(n499) );
  NOR2BX1TS U563 ( .AN(n596), .B(n643), .Y(n496) );
  AOI31XLTS U564 ( .A0(n318), .A1(n499), .A2(n496), .B0(reset), .Y(rf_raa[1])
         );
  OR2X1TS U565 ( .A(n319), .B(rf_raa[1]), .Y(rf_raa[5]) );
  CLKBUFX2TS U566 ( .A(rf_raa[5]), .Y(rf_rea) );
  AOI31XLTS U567 ( .A0(n580), .A1(n321), .A2(start), .B0(n320), .Y(n324) );
  AOI31XLTS U568 ( .A0(mode[1]), .A1(n641), .A2(n639), .B0(n322), .Y(n323) );
  NOR4BXLTS U569 ( .AN(n324), .B(n553), .C(n460), .D(n323), .Y(n325) );
  OAI211XLTS U570 ( .A0(comp2_g), .A1(n326), .B0(n325), .C0(n464), .Y(n327) );
  AOI211XLTS U571 ( .A0(N2139), .A1(n328), .B0(n477), .C0(n327), .Y(n351) );
  INVX2TS U572 ( .A(sumor), .Y(n329) );
  AOI22X1TS U573 ( .A0(comp1_g), .A1(n331), .B0(n330), .B1(n329), .Y(n339) );
  NAND3XLTS U574 ( .A(n334), .B(n333), .C(n332), .Y(n337) );
  INVX2TS U575 ( .A(n335), .Y(n607) );
  AOI211XLTS U576 ( .A0(mq47), .A1(n337), .B0(n336), .C0(n607), .Y(n338) );
  OAI211XLTS U577 ( .A0(st), .A1(n480), .B0(n339), .C0(n338), .Y(n349) );
  OAI211XLTS U578 ( .A0(mq47), .A1(n340), .B0(n597), .C0(n613), .Y(n341) );
  AOI211XLTS U579 ( .A0(n344), .A1(n343), .B0(n342), .C0(n341), .Y(n345) );
  NAND3XLTS U580 ( .A(n347), .B(n346), .C(n345), .Y(n348) );
  AOI211XLTS U581 ( .A0(n360), .A1(n462), .B0(n349), .C0(n348), .Y(n350) );
  AOI31XLTS U582 ( .A0(n352), .A1(n351), .A2(n350), .B0(reset), .Y(N2445) );
  AOI211XLTS U583 ( .A0(N2131), .A1(n355), .B0(n354), .C0(n353), .Y(n386) );
  AOI22X1TS U584 ( .A0(mq47), .A1(n356), .B0(n473), .B1(msb), .Y(n358) );
  OAI211XLTS U585 ( .A0(n359), .A1(n638), .B0(n358), .C0(n357), .Y(n380) );
  AOI22X1TS U586 ( .A0(n631), .A1(n362), .B0(n361), .B1(n360), .Y(n378) );
  INVX2TS U587 ( .A(r31), .Y(n365) );
  AOI22X1TS U588 ( .A0(n366), .A1(n365), .B0(n364), .B1(n363), .Y(n377) );
  AOI32X1TS U589 ( .A0(n439), .A1(n599), .A2(n367), .B0(n408), .B1(n599), .Y(
        n368) );
  NOR4XLTS U590 ( .A(n460), .B(n448), .C(n369), .D(n368), .Y(n376) );
  INVX2TS U591 ( .A(n370), .Y(n374) );
  AOI21X1TS U592 ( .A0(n371), .A1(n610), .B0(n383), .Y(n373) );
  AOI211XLTS U593 ( .A0(N2152), .A1(n374), .B0(n373), .C0(n372), .Y(n375) );
  NAND4XLTS U594 ( .A(n378), .B(n377), .C(n376), .D(n375), .Y(n379) );
  NOR4BXLTS U595 ( .AN(n382), .B(n381), .C(n380), .D(n379), .Y(n385) );
  OAI2BB1X1TS U596 ( .A0N(n620), .A1N(n611), .B0(n383), .Y(n384) );
  AOI31XLTS U597 ( .A0(n386), .A1(n385), .A2(n384), .B0(reset), .Y(N2447) );
  OAI32X1TS U598 ( .A0(reset), .A1(state[1]), .A2(n387), .B0(n568), .B1(reset), 
        .Y(n388) );
  CLKBUFX2TS U599 ( .A(n388), .Y(reg_ma) );
  INVX2TS U600 ( .A(reg_ma), .Y(n541) );
  INVX2TS U601 ( .A(n541), .Y(mux15) );
  INVX2TS U602 ( .A(n541), .Y(reg_sa) );
  CLKAND2X2TS U603 ( .A(n557), .B(state[4]), .Y(n447) );
  AOI222XLTS U604 ( .A0(n579), .A1(n447), .B0(n578), .B1(n571), .C0(n401), 
        .C1(n530), .Y(n390) );
  AOI221XLTS U605 ( .A0(state[8]), .A1(n391), .B0(n397), .B1(n390), .C0(n590), 
        .Y(n392) );
  AOI31XLTS U606 ( .A0(n417), .A1(n415), .A2(n393), .B0(n392), .Y(n404) );
  OAI2BB2XLTS U607 ( .B0(n469), .B1(n394), .A0N(n578), .A1N(n393), .Y(n398) );
  OAI21XLTS U608 ( .A0(n513), .A1(n397), .B0(n484), .Y(n395) );
  AOI222XLTS U609 ( .A0(n398), .A1(n397), .B0(n396), .B1(n571), .C0(n395), 
        .C1(n401), .Y(n399) );
  OAI21XLTS U610 ( .A0(n399), .A1(n590), .B0(state[3]), .Y(n400) );
  AOI31XLTS U611 ( .A0(n417), .A1(n402), .A2(n401), .B0(n400), .Y(n403) );
  AOI211XLTS U612 ( .A0(n404), .A1(n416), .B0(reset), .C0(n403), .Y(n405) );
  CLKBUFX2TS U613 ( .A(n405), .Y(reg_currterm) );
  INVX2TS U614 ( .A(reg_mc), .Y(n542) );
  INVX2TS U615 ( .A(n542), .Y(reg_sc) );
  OAI22X1TS U616 ( .A0(n584), .A1(n408), .B0(n556), .B1(n407), .Y(n414) );
  NOR3XLTS U617 ( .A(n411), .B(n410), .C(n409), .Y(n413) );
  AOI211XLTS U618 ( .A0(n415), .A1(n414), .B0(n413), .C0(n412), .Y(n420) );
  OAI31X1TS U619 ( .A0(n417), .A1(n416), .A2(n446), .B0(n445), .Y(n418) );
  NOR2XLTS U620 ( .A(n563), .B(n561), .Y(n583) );
  AOI32X1TS U621 ( .A0(n571), .A1(n422), .A2(n418), .B0(n583), .B1(n422), .Y(
        n419) );
  NAND4XLTS U622 ( .A(n420), .B(n442), .C(n598), .D(n419), .Y(n421) );
  INVX2TS U623 ( .A(n489), .Y(n425) );
  NAND2X1TS U624 ( .A(n531), .B(n530), .Y(n423) );
  NAND2X1TS U625 ( .A(n569), .B(n422), .Y(n498) );
  AOI32X1TS U626 ( .A0(n593), .A1(n423), .A2(n498), .B0(n525), .B1(n423), .Y(
        n424) );
  AOI32X1TS U627 ( .A0(n524), .A1(state[5]), .A2(n434), .B0(n424), .B1(n559), 
        .Y(n485) );
  OAI32X1TS U628 ( .A0(reset), .A1(n425), .A2(n485), .B0(n499), .B1(reset), 
        .Y(rf_rab_5) );
  CLKBUFX2TS U629 ( .A(rf_rab_5), .Y(reg_mb) );
  INVX2TS U630 ( .A(reg_mb), .Y(n543) );
  INVX2TS U631 ( .A(n543), .Y(reg_sb) );
  INVX2TS U632 ( .A(n426), .Y(n551) );
  NOR2XLTS U633 ( .A(reset), .B(n551), .Y(n427) );
  CLKBUFX2TS U634 ( .A(n427), .Y(reg_numbit) );
  NAND2X1TS U635 ( .A(n471), .B(n430), .Y(n433) );
  INVX2TS U636 ( .A(n433), .Y(mux4[1]) );
  INVX2TS U637 ( .A(n433), .Y(mux5) );
  NAND3XLTS U638 ( .A(n433), .B(n432), .C(n431), .Y(sr_mt[0]) );
  NAND2X1TS U639 ( .A(n435), .B(n434), .Y(n437) );
  AOI31XLTS U640 ( .A0(n438), .A1(n437), .A2(n436), .B0(reset), .Y(mux10) );
  OAI21XLTS U641 ( .A0(n439), .A1(n527), .B0(n442), .Y(n440) );
  AOI211XLTS U642 ( .A0(n471), .A1(n440), .B0(mux2[0]), .C0(mux21[0]), .Y(n441) );
  NAND2X1TS U643 ( .A(n601), .B(n441), .Y(mux2[1]) );
  AOI21X1TS U644 ( .A0(n495), .A1(n442), .B0(reset), .Y(mux2[2]) );
  NOR2XLTS U645 ( .A(reset), .B(n443), .Y(mux23) );
  OAI33XLTS U646 ( .A0(state[6]), .A1(n563), .A2(n556), .B0(n536), .B1(n528), 
        .B2(state[7]), .Y(n444) );
  NAND2X1TS U647 ( .A(state[5]), .B(n444), .Y(n570) );
  OAI21XLTS U648 ( .A0(n446), .A1(n528), .B0(n445), .Y(n581) );
  OAI2BB2XLTS U649 ( .B0(n508), .B1(n570), .A0N(n447), .A1N(n581), .Y(n450) );
  AOI211XLTS U650 ( .A0(state[1]), .A1(n450), .B0(n449), .C0(n448), .Y(n451)
         );
  NOR2XLTS U651 ( .A(reset), .B(n451), .Y(mux3[2]) );
  CLKAND2X2TS U652 ( .A(n452), .B(n471), .Y(rf_wa[0]) );
  OR2X1TS U653 ( .A(rf_wa[0]), .B(rf_wa[1]), .Y(rf_wa_5) );
  INVX2TS U654 ( .A(n455), .Y(n453) );
  AOI21X1TS U655 ( .A0(n659), .A1(n453), .B0(reset), .Y(mux17_0) );
  AOI31X1TS U656 ( .A0(n458), .A1(n457), .A2(n456), .B0(reset), .Y(alu2[1]) );
  OR2X1TS U657 ( .A(mux17[2]), .B(alu2[1]), .Y(alu2[2]) );
  OAI21XLTS U658 ( .A0(n553), .A1(n459), .B0(n471), .Y(n609) );
  INVX2TS U659 ( .A(mux21[0]), .Y(n594) );
  NAND3XLTS U660 ( .A(n609), .B(n594), .C(n595), .Y(sr_res[0]) );
  AOI2BB1XLTS U661 ( .A0N(n461), .A1N(n460), .B0(reset), .Y(sr_res[1]) );
  AOI21X1TS U662 ( .A0(n475), .A1(n502), .B0(reset), .Y(mux9[2]) );
  OAI31X1TS U663 ( .A0(n462), .A1(mux9[2]), .A2(n473), .B0(n471), .Y(n463) );
  INVX2TS U664 ( .A(ssr_ms0[1]), .Y(n472) );
  NAND2X1TS U665 ( .A(n463), .B(n472), .Y(reg_es0) );
  CLKAND2X2TS U666 ( .A(n465), .B(n464), .Y(n467) );
  NOR2BX1TS U667 ( .AN(n474), .B(n466), .Y(n548) );
  AOI31XLTS U668 ( .A0(n475), .A1(n467), .A2(n548), .B0(reset), .Y(mux9[0]) );
  NAND3XLTS U669 ( .A(n489), .B(state[2]), .C(n535), .Y(n468) );
  OAI21XLTS U670 ( .A0(n469), .A1(n570), .B0(n468), .Y(n470) );
  NAND3XLTS U671 ( .A(state[1]), .B(n471), .C(n470), .Y(n575) );
  OAI21XLTS U672 ( .A0(reset), .A1(n502), .B0(n575), .Y(mux6[1]) );
  NAND3BXLTS U673 ( .AN(mux6[1]), .B(n609), .C(n472), .Y(alu1[0]) );
  INVX2TS U674 ( .A(n473), .Y(n550) );
  AOI31X1TS U675 ( .A0(n551), .A1(n480), .A2(n479), .B0(reset), .Y(alu1[1]) );
  OR2X1TS U676 ( .A(mux6[1]), .B(alu1[1]), .Y(alu1[2]) );
  AOI32X1TS U677 ( .A0(n571), .A1(n482), .A2(n524), .B0(n481), .B1(n482), .Y(
        n493) );
  OAI22X1TS U678 ( .A0(n556), .A1(n484), .B0(n483), .B1(n508), .Y(n488) );
  OAI31X1TS U679 ( .A0(state[2]), .A1(state[1]), .A2(n486), .B0(n485), .Y(n487) );
  AOI32X1TS U680 ( .A0(state[5]), .A1(n489), .A2(n488), .B0(n487), .B1(n489), 
        .Y(n492) );
  OAI221XLTS U681 ( .A0(state[1]), .A1(n498), .B0(n590), .B1(n569), .C0(n490), 
        .Y(n491) );
  AOI31XLTS U682 ( .A0(n493), .A1(n492), .A2(n491), .B0(reset), .Y(rf_reb) );
  AOI21X1TS U683 ( .A0(n495), .A1(n494), .B0(reset), .Y(rf_raa[0]) );
  OAI32X1TS U684 ( .A0(reset), .A1(n498), .A2(n497), .B0(n496), .B1(reset), 
        .Y(rf_rab[1]) );
  NOR2XLTS U685 ( .A(reset), .B(n499), .Y(rf_rab[0]) );
  AOI22X1TS U686 ( .A0(n501), .A1(state[4]), .B0(n500), .B1(n569), .Y(n521) );
  INVX2TS U687 ( .A(n502), .Y(n616) );
  OAI22X1TS U688 ( .A0(n505), .A1(n508), .B0(n504), .B1(n503), .Y(n506) );
  AOI211XLTS U689 ( .A0(n628), .A1(state[4]), .B0(n616), .C0(n506), .Y(n520)
         );
  AOI22X1TS U690 ( .A0(state[6]), .A1(n507), .B0(n514), .B1(n536), .Y(n512) );
  OAI21XLTS U691 ( .A0(n631), .A1(n590), .B0(n508), .Y(n510) );
  AOI211XLTS U692 ( .A0(n569), .A1(n590), .B0(state[4]), .C0(n584), .Y(n509)
         );
  AOI32X1TS U693 ( .A0(n515), .A1(n536), .A2(n510), .B0(state[6]), .B1(n509), 
        .Y(n511) );
  OAI31X1TS U694 ( .A0(state[1]), .A1(n513), .A2(n512), .B0(n511), .Y(n518) );
  AOI22X1TS U695 ( .A0(n515), .A1(n571), .B0(n514), .B1(n569), .Y(n516) );
  OAI31X1TS U696 ( .A0(n516), .A1(n536), .A2(n590), .B0(state[5]), .Y(n517) );
  OAI211XLTS U697 ( .A0(state[5]), .A1(n518), .B0(n563), .C0(n517), .Y(n519)
         );
  AOI31XLTS U698 ( .A0(n521), .A1(n520), .A2(n519), .B0(reset), .Y(reg_ss0) );
  AOI211XLTS U699 ( .A0(state[2]), .A1(state[1]), .B0(state[0]), .C0(n563), 
        .Y(n537) );
  AOI22X1TS U700 ( .A0(n631), .A1(n524), .B0(n580), .B1(n523), .Y(n533) );
  OAI22X1TS U701 ( .A0(n528), .A1(n527), .B0(n526), .B1(n525), .Y(n529) );
  AOI21X1TS U702 ( .A0(n531), .A1(n530), .B0(n529), .Y(n532) );
  AOI221XLTS U703 ( .A0(state[5]), .A1(n533), .B0(n559), .B1(n532), .C0(
        state[7]), .Y(n534) );
  AOI32X1TS U704 ( .A0(n537), .A1(n536), .A2(n535), .B0(n534), .B1(n536), .Y(
        n538) );
  AOI31X1TS U705 ( .A0(n540), .A1(n539), .A2(n538), .B0(reset), .Y(reg_index)
         );
  INVX2TS U706 ( .A(n541), .Y(reg_ea) );
  INVX2TS U707 ( .A(n433), .Y(reg_st) );
  INVX2TS U708 ( .A(n433), .Y(reg_ss) );
  INVX2TS U709 ( .A(n542), .Y(reg_ec) );
  INVX2TS U710 ( .A(n543), .Y(reg_eb) );
  NOR2XLTS U711 ( .A(n545), .B(n544), .Y(n547) );
  OAI21XLTS U712 ( .A0(reset), .A1(n547), .B0(n601), .Y(mux13[1]) );
  AOI31XLTS U713 ( .A0(n596), .A1(n547), .A2(n546), .B0(reset), .Y(mux13[2])
         );
  AOI31XLTS U714 ( .A0(n549), .A1(n548), .A2(n550), .B0(reset), .Y(mux8[0]) );
  AOI21X1TS U715 ( .A0(n551), .A1(n550), .B0(reset), .Y(mux9[1]) );
  INVX2TS U716 ( .A(n433), .Y(reg_es) );
  INVX2TS U717 ( .A(n433), .Y(reg_et) );
  NOR2XLTS U718 ( .A(n552), .B(reset), .Y(counterii[2]) );
  OR2X1TS U719 ( .A(sr_mq[0]), .B(sr_mp[0]), .Y(alu2[0]) );
  AOI21X1TS U720 ( .A0(n629), .A1(n554), .B0(n553), .Y(n567) );
  OAI22X1TS U721 ( .A0(n557), .A1(n556), .B0(n584), .B1(n555), .Y(n558) );
  AOI32X1TS U722 ( .A0(n560), .A1(state[5]), .A2(n577), .B0(n559), .B1(n558), 
        .Y(n562) );
  OAI32X1TS U723 ( .A0(state[1]), .A1(state[6]), .A2(n562), .B0(n561), .B1(
        state[1]), .Y(n564) );
  AOI22X1TS U724 ( .A0(n565), .A1(n571), .B0(n564), .B1(n563), .Y(n566) );
  AOI31XLTS U725 ( .A0(n568), .A1(n567), .A2(n566), .B0(reset), .Y(mux19) );
  OAI2BB2XLTS U726 ( .B0(n631), .B1(n570), .A0N(n569), .A1N(n581), .Y(n574) );
  AOI222XLTS U727 ( .A0(n574), .A1(n590), .B0(n629), .B1(n573), .C0(n572), 
        .C1(n571), .Y(n576) );
  OAI21XLTS U728 ( .A0(reset), .A1(n576), .B0(n575), .Y(mux12[1]) );
  AOI22X1TS U729 ( .A0(n580), .A1(n579), .B0(n578), .B1(n577), .Y(n587) );
  AOI22X1TS U730 ( .A0(state[0]), .A1(n583), .B0(n582), .B1(n581), .Y(n586) );
  AOI32X1TS U731 ( .A0(n587), .A1(n586), .A2(n585), .B0(n584), .B1(n586), .Y(
        n589) );
  AOI211XLTS U732 ( .A0(n590), .A1(n589), .B0(n616), .C0(n588), .Y(n591) );
  OAI32X1TS U733 ( .A0(reset), .A1(n593), .A2(n592), .B0(n591), .B1(reset), 
        .Y(mux11) );
  CLKAND2X2TS U734 ( .A(n598), .B(n597), .Y(n600) );
  AOI31XLTS U735 ( .A0(n600), .A1(n599), .A2(n602), .B0(reset), .Y(mux14[0])
         );
  NAND2X1TS U736 ( .A(n602), .B(n601), .Y(reg_i) );
  NOR2XLTS U737 ( .A(n604), .B(n603), .Y(n605) );
  AOI21X1TS U738 ( .A0(n606), .A1(n605), .B0(reset), .Y(mux6[0]) );
  AOI2BB1XLTS U739 ( .A0N(n607), .A1N(n642), .B0(reset), .Y(reg_e) );
  NAND2X1TS U740 ( .A(n609), .B(n608), .Y(mux8[2]) );
  OAI22X1TS U741 ( .A0(n612), .A1(n611), .B0(n610), .B1(n644), .Y(n622) );
  INVX2TS U742 ( .A(n613), .Y(n615) );
  AOI211XLTS U743 ( .A0(ms0_23), .A1(n616), .B0(n615), .C0(n614), .Y(n617) );
  OAI211XLTS U744 ( .A0(n620), .A1(n619), .B0(n618), .C0(n617), .Y(n621) );
  NOR4BXLTS U745 ( .AN(n624), .B(n623), .C(n622), .D(n621), .Y(n655) );
  AOI22X1TS U746 ( .A0(n631), .A1(n627), .B0(n626), .B1(n625), .Y(n633) );
  AOI22X1TS U747 ( .A0(n631), .A1(n630), .B0(n629), .B1(n628), .Y(n632) );
  OAI211XLTS U748 ( .A0(n635), .A1(n634), .B0(n633), .C0(n632), .Y(n652) );
  OAI211XLTS U749 ( .A0(mode[0]), .A1(n640), .B0(n637), .C0(n636), .Y(n651) );
  OA22X1TS U750 ( .A0(n641), .A1(n640), .B0(n639), .B1(n638), .Y(n647) );
  AOI211XLTS U751 ( .A0(n645), .A1(n644), .B0(n643), .C0(n642), .Y(n646) );
  OAI211XLTS U752 ( .A0(n649), .A1(n648), .B0(n647), .C0(n646), .Y(n650) );
  NOR4XLTS U753 ( .A(n653), .B(n652), .C(n651), .D(n650), .Y(n654) );
  AOI21X1TS U754 ( .A0(n655), .A1(n654), .B0(reset), .Y(N2448) );
  NAND4XLTS U755 ( .A(n659), .B(n658), .C(n657), .D(n656), .Y(N2444) );
endmodule


module mult32_1 ( A, B, Product );
  input [31:0] A;
  input [31:0] B;
  output [63:0] Product;
  wire   \mult_x_1/n1250 , \mult_x_1/n1249 , \mult_x_1/n1248 ,
         \mult_x_1/n1247 , \mult_x_1/n1246 , \mult_x_1/n1245 ,
         \mult_x_1/n1244 , \mult_x_1/n1243 , \mult_x_1/n1242 ,
         \mult_x_1/n1241 , \mult_x_1/n1240 , \mult_x_1/n1239 ,
         \mult_x_1/n1238 , \mult_x_1/n1237 , \mult_x_1/n1236 ,
         \mult_x_1/n1235 , \mult_x_1/n1234 , \mult_x_1/n1233 ,
         \mult_x_1/n1232 , \mult_x_1/n1231 , \mult_x_1/n1218 ,
         \mult_x_1/n1217 , \mult_x_1/n1216 , \mult_x_1/n1215 ,
         \mult_x_1/n1214 , \mult_x_1/n1213 , \mult_x_1/n1212 ,
         \mult_x_1/n1211 , \mult_x_1/n1210 , \mult_x_1/n1209 ,
         \mult_x_1/n1208 , \mult_x_1/n1207 , \mult_x_1/n1206 ,
         \mult_x_1/n1205 , \mult_x_1/n1204 , \mult_x_1/n1203 ,
         \mult_x_1/n1202 , \mult_x_1/n1201 , \mult_x_1/n1200 ,
         \mult_x_1/n1199 , \mult_x_1/n1198 , \mult_x_1/n1197 ,
         \mult_x_1/n1196 , \mult_x_1/n1180 , \mult_x_1/n1179 ,
         \mult_x_1/n1178 , \mult_x_1/n1177 , \mult_x_1/n1176 ,
         \mult_x_1/n1175 , \mult_x_1/n1174 , \mult_x_1/n1173 ,
         \mult_x_1/n1172 , \mult_x_1/n1171 , \mult_x_1/n1170 ,
         \mult_x_1/n1169 , \mult_x_1/n1168 , \mult_x_1/n1167 ,
         \mult_x_1/n1166 , \mult_x_1/n1165 , \mult_x_1/n1164 ,
         \mult_x_1/n1163 , \mult_x_1/n1162 , \mult_x_1/n1161 ,
         \mult_x_1/n1148 , \mult_x_1/n1147 , \mult_x_1/n1146 ,
         \mult_x_1/n1145 , \mult_x_1/n1144 , \mult_x_1/n1143 ,
         \mult_x_1/n1142 , \mult_x_1/n1141 , \mult_x_1/n1140 ,
         \mult_x_1/n1139 , \mult_x_1/n1138 , \mult_x_1/n1137 ,
         \mult_x_1/n1136 , \mult_x_1/n1135 , \mult_x_1/n1134 ,
         \mult_x_1/n1133 , \mult_x_1/n1132 , \mult_x_1/n1131 ,
         \mult_x_1/n1130 , \mult_x_1/n1129 , \mult_x_1/n1128 ,
         \mult_x_1/n1127 , \mult_x_1/n1126 , \mult_x_1/n1110 ,
         \mult_x_1/n1109 , \mult_x_1/n1108 , \mult_x_1/n1107 ,
         \mult_x_1/n1106 , \mult_x_1/n1105 , \mult_x_1/n1104 ,
         \mult_x_1/n1103 , \mult_x_1/n1102 , \mult_x_1/n1101 ,
         \mult_x_1/n1100 , \mult_x_1/n1099 , \mult_x_1/n1098 ,
         \mult_x_1/n1097 , \mult_x_1/n1096 , \mult_x_1/n1095 ,
         \mult_x_1/n1094 , \mult_x_1/n1093 , \mult_x_1/n1092 ,
         \mult_x_1/n1091 , \mult_x_1/n1078 , \mult_x_1/n1077 ,
         \mult_x_1/n1076 , \mult_x_1/n1075 , \mult_x_1/n1074 ,
         \mult_x_1/n1073 , \mult_x_1/n1072 , \mult_x_1/n1071 ,
         \mult_x_1/n1070 , \mult_x_1/n1069 , \mult_x_1/n1068 ,
         \mult_x_1/n1067 , \mult_x_1/n1066 , \mult_x_1/n1065 ,
         \mult_x_1/n1064 , \mult_x_1/n1063 , \mult_x_1/n1062 ,
         \mult_x_1/n1061 , \mult_x_1/n1060 , \mult_x_1/n1059 ,
         \mult_x_1/n1058 , \mult_x_1/n1057 , \mult_x_1/n1056 ,
         \mult_x_1/n1032 , \mult_x_1/n1031 , \mult_x_1/n1030 ,
         \mult_x_1/n1029 , \mult_x_1/n1028 , \mult_x_1/n1027 ,
         \mult_x_1/n1025 , \mult_x_1/n1024 , \mult_x_1/n1023 ,
         \mult_x_1/n1022 , \mult_x_1/n1021 , \mult_x_1/n798 , \mult_x_1/n796 ,
         \mult_x_1/n795 , \mult_x_1/n793 , \mult_x_1/n792 , \mult_x_1/n791 ,
         \mult_x_1/n790 , \mult_x_1/n788 , \mult_x_1/n787 , \mult_x_1/n786 ,
         \mult_x_1/n785 , \mult_x_1/n783 , \mult_x_1/n782 , \mult_x_1/n781 ,
         \mult_x_1/n778 , \mult_x_1/n776 , \mult_x_1/n775 , \mult_x_1/n774 ,
         \mult_x_1/n771 , \mult_x_1/n769 , \mult_x_1/n768 , \mult_x_1/n767 ,
         \mult_x_1/n765 , \mult_x_1/n764 , \mult_x_1/n763 , \mult_x_1/n762 ,
         \mult_x_1/n761 , \mult_x_1/n760 , \mult_x_1/n759 , \mult_x_1/n757 ,
         \mult_x_1/n756 , \mult_x_1/n755 , \mult_x_1/n754 , \mult_x_1/n753 ,
         \mult_x_1/n752 , \mult_x_1/n751 , \mult_x_1/n749 , \mult_x_1/n748 ,
         \mult_x_1/n747 , \mult_x_1/n746 , \mult_x_1/n745 , \mult_x_1/n744 ,
         \mult_x_1/n743 , \mult_x_1/n741 , \mult_x_1/n740 , \mult_x_1/n739 ,
         \mult_x_1/n738 , \mult_x_1/n737 , \mult_x_1/n736 , \mult_x_1/n733 ,
         \mult_x_1/n731 , \mult_x_1/n730 , \mult_x_1/n729 , \mult_x_1/n728 ,
         \mult_x_1/n727 , \mult_x_1/n726 , \mult_x_1/n723 , \mult_x_1/n721 ,
         \mult_x_1/n720 , \mult_x_1/n719 , \mult_x_1/n718 , \mult_x_1/n717 ,
         \mult_x_1/n716 , \mult_x_1/n714 , \mult_x_1/n713 , \mult_x_1/n712 ,
         \mult_x_1/n711 , \mult_x_1/n710 , \mult_x_1/n709 , \mult_x_1/n708 ,
         \mult_x_1/n707 , \mult_x_1/n706 , \mult_x_1/n705 , \mult_x_1/n703 ,
         \mult_x_1/n702 , \mult_x_1/n701 , \mult_x_1/n700 , \mult_x_1/n699 ,
         \mult_x_1/n698 , \mult_x_1/n697 , \mult_x_1/n696 , \mult_x_1/n695 ,
         \mult_x_1/n694 , \mult_x_1/n692 , \mult_x_1/n691 , \mult_x_1/n690 ,
         \mult_x_1/n689 , \mult_x_1/n688 , \mult_x_1/n687 , \mult_x_1/n686 ,
         \mult_x_1/n685 , \mult_x_1/n684 , \mult_x_1/n683 , \mult_x_1/n681 ,
         \mult_x_1/n680 , \mult_x_1/n679 , \mult_x_1/n678 , \mult_x_1/n677 ,
         \mult_x_1/n676 , \mult_x_1/n675 , \mult_x_1/n674 , \mult_x_1/n673 ,
         \mult_x_1/n670 , \mult_x_1/n668 , \mult_x_1/n667 , \mult_x_1/n666 ,
         \mult_x_1/n665 , \mult_x_1/n664 , \mult_x_1/n663 , \mult_x_1/n662 ,
         \mult_x_1/n661 , \mult_x_1/n660 , \mult_x_1/n657 , \mult_x_1/n655 ,
         \mult_x_1/n654 , \mult_x_1/n653 , \mult_x_1/n652 , \mult_x_1/n651 ,
         \mult_x_1/n650 , \mult_x_1/n649 , \mult_x_1/n648 , \mult_x_1/n647 ,
         \mult_x_1/n644 , \mult_x_1/n642 , \mult_x_1/n641 , \mult_x_1/n640 ,
         \mult_x_1/n639 , \mult_x_1/n638 , \mult_x_1/n637 , \mult_x_1/n636 ,
         \mult_x_1/n635 , \mult_x_1/n634 , \mult_x_1/n631 , \mult_x_1/n628 ,
         \mult_x_1/n627 , \mult_x_1/n626 , \mult_x_1/n625 , \mult_x_1/n624 ,
         \mult_x_1/n623 , \mult_x_1/n622 , \mult_x_1/n621 , \mult_x_1/n620 ,
         \mult_x_1/n617 , \mult_x_1/n614 , \mult_x_1/n613 , \mult_x_1/n612 ,
         \mult_x_1/n611 , \mult_x_1/n610 , \mult_x_1/n609 , \mult_x_1/n608 ,
         \mult_x_1/n607 , \mult_x_1/n606 , \mult_x_1/n603 , \mult_x_1/n600 ,
         \mult_x_1/n599 , \mult_x_1/n598 , \mult_x_1/n597 , \mult_x_1/n596 ,
         \mult_x_1/n595 , \mult_x_1/n594 , \mult_x_1/n593 , \mult_x_1/n592 ,
         \mult_x_1/n589 , \mult_x_1/n586 , \mult_x_1/n585 , \mult_x_1/n584 ,
         \mult_x_1/n583 , \mult_x_1/n582 , \mult_x_1/n581 , \mult_x_1/n580 ,
         \mult_x_1/n579 , \mult_x_1/n578 , \mult_x_1/n575 , \mult_x_1/n572 ,
         \mult_x_1/n571 , \mult_x_1/n570 , \mult_x_1/n569 , \mult_x_1/n568 ,
         \mult_x_1/n567 , \mult_x_1/n566 , \mult_x_1/n565 , \mult_x_1/n564 ,
         \mult_x_1/n561 , \mult_x_1/n558 , \mult_x_1/n557 , \mult_x_1/n556 ,
         \mult_x_1/n555 , \mult_x_1/n554 , \mult_x_1/n553 , \mult_x_1/n552 ,
         \mult_x_1/n551 , \mult_x_1/n550 , \mult_x_1/n547 , \mult_x_1/n546 ,
         \mult_x_1/n544 , \mult_x_1/n543 , \mult_x_1/n542 , \mult_x_1/n541 ,
         \mult_x_1/n540 , \mult_x_1/n539 , \mult_x_1/n538 , \mult_x_1/n537 ,
         \mult_x_1/n536 , \mult_x_1/n533 , \mult_x_1/n530 , \mult_x_1/n529 ,
         \mult_x_1/n528 , \mult_x_1/n527 , \mult_x_1/n526 , \mult_x_1/n525 ,
         \mult_x_1/n524 , \mult_x_1/n523 , \mult_x_1/n522 , \mult_x_1/n519 ,
         \mult_x_1/n516 , \mult_x_1/n515 , \mult_x_1/n514 , \mult_x_1/n513 ,
         \mult_x_1/n512 , \mult_x_1/n511 , \mult_x_1/n510 , \mult_x_1/n509 ,
         \mult_x_1/n508 , \mult_x_1/n505 , \mult_x_1/n502 , \mult_x_1/n501 ,
         \mult_x_1/n500 , \mult_x_1/n499 , \mult_x_1/n498 , \mult_x_1/n497 ,
         \mult_x_1/n496 , \mult_x_1/n495 , \mult_x_1/n494 , \mult_x_1/n491 ,
         \mult_x_1/n488 , \mult_x_1/n487 , \mult_x_1/n486 , \mult_x_1/n485 ,
         \mult_x_1/n484 , \mult_x_1/n483 , \mult_x_1/n482 , \mult_x_1/n481 ,
         \mult_x_1/n480 , \mult_x_1/n475 , \mult_x_1/n474 , \mult_x_1/n473 ,
         \mult_x_1/n472 , \mult_x_1/n471 , \mult_x_1/n470 , \mult_x_1/n469 ,
         \mult_x_1/n468 , \mult_x_1/n467 , \mult_x_1/n464 , \mult_x_1/n463 ,
         \mult_x_1/n461 , \mult_x_1/n460 , \mult_x_1/n459 , \mult_x_1/n458 ,
         \mult_x_1/n457 , \mult_x_1/n456 , \mult_x_1/n455 , \mult_x_1/n454 ,
         \mult_x_1/n453 , \mult_x_1/n452 , \mult_x_1/n450 , \mult_x_1/n449 ,
         \mult_x_1/n448 , \mult_x_1/n447 , \mult_x_1/n446 , \mult_x_1/n445 ,
         \mult_x_1/n444 , \mult_x_1/n443 , \mult_x_1/n442 , \mult_x_1/n438 ,
         \mult_x_1/n435 , \mult_x_1/n434 , \mult_x_1/n433 , \mult_x_1/n432 ,
         \mult_x_1/n431 , \mult_x_1/n430 , \mult_x_1/n425 , \mult_x_1/n424 ,
         \mult_x_1/n422 , \mult_x_1/n421 , \mult_x_1/n420 , \mult_x_1/n419 ,
         \mult_x_1/n418 , \mult_x_1/n417 , \mult_x_1/n414 , \mult_x_1/n413 ,
         \mult_x_1/n411 , \mult_x_1/n410 , \mult_x_1/n409 , \mult_x_1/n408 ,
         \mult_x_1/n407 , \mult_x_1/n406 , \mult_x_1/n404 , \mult_x_1/n401 ,
         \mult_x_1/n400 , \mult_x_1/n399 , \mult_x_1/n398 , \mult_x_1/n397 ,
         \mult_x_1/n396 , \mult_x_1/n390 , \mult_x_1/n389 , \mult_x_1/n388 ,
         \mult_x_1/n387 , \mult_x_1/n386 , \mult_x_1/n385 , \mult_x_1/n382 ,
         \mult_x_1/n381 , \mult_x_1/n379 , \mult_x_1/n378 , \mult_x_1/n377 ,
         \mult_x_1/n373 , \mult_x_1/n370 , \mult_x_1/n369 , \mult_x_1/n368 ,
         \mult_x_1/n363 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1034, n1035, n1036;

  CMPR42X1TS \mult_x_1/U485  ( .A(\mult_x_1/n795 ), .B(\mult_x_1/n1218 ), .C(
        \mult_x_1/n798 ), .D(\mult_x_1/n1250 ), .ICI(\mult_x_1/n796 ), .S(
        \mult_x_1/n793 ), .ICO(\mult_x_1/n791 ), .CO(\mult_x_1/n792 ) );
  CMPR42X1TS \mult_x_1/U483  ( .A(\mult_x_1/n790 ), .B(\mult_x_1/n1217 ), .C(
        \mult_x_1/n791 ), .D(\mult_x_1/n1249 ), .ICI(\mult_x_1/n792 ), .S(
        \mult_x_1/n788 ), .ICO(\mult_x_1/n786 ), .CO(\mult_x_1/n787 ) );
  CMPR42X1TS \mult_x_1/U481  ( .A(\mult_x_1/n785 ), .B(\mult_x_1/n1216 ), .C(
        \mult_x_1/n786 ), .D(\mult_x_1/n1248 ), .ICI(\mult_x_1/n787 ), .S(
        \mult_x_1/n783 ), .ICO(\mult_x_1/n781 ), .CO(\mult_x_1/n782 ) );
  CMPR42X1TS \mult_x_1/U478  ( .A(\mult_x_1/n778 ), .B(\mult_x_1/n781 ), .C(
        \mult_x_1/n1215 ), .D(\mult_x_1/n1247 ), .ICI(\mult_x_1/n782 ), .S(
        \mult_x_1/n776 ), .ICO(\mult_x_1/n774 ), .CO(\mult_x_1/n775 ) );
  CMPR42X1TS \mult_x_1/U475  ( .A(\mult_x_1/n771 ), .B(\mult_x_1/n774 ), .C(
        \mult_x_1/n1214 ), .D(\mult_x_1/n1246 ), .ICI(\mult_x_1/n775 ), .S(
        \mult_x_1/n769 ), .ICO(\mult_x_1/n767 ), .CO(\mult_x_1/n768 ) );
  CMPR42X1TS \mult_x_1/U472  ( .A(\mult_x_1/n764 ), .B(\mult_x_1/n767 ), .C(
        \mult_x_1/n1213 ), .D(\mult_x_1/n1245 ), .ICI(\mult_x_1/n768 ), .S(
        \mult_x_1/n762 ), .ICO(\mult_x_1/n760 ), .CO(\mult_x_1/n761 ) );
  CMPR42X1TS \mult_x_1/U470  ( .A(\mult_x_1/n759 ), .B(\mult_x_1/n1148 ), .C(
        \mult_x_1/n765 ), .D(\mult_x_1/n1180 ), .ICI(\mult_x_1/n763 ), .S(
        \mult_x_1/n757 ), .ICO(\mult_x_1/n755 ), .CO(\mult_x_1/n756 ) );
  CMPR42X1TS \mult_x_1/U469  ( .A(\mult_x_1/n757 ), .B(\mult_x_1/n760 ), .C(
        \mult_x_1/n1212 ), .D(\mult_x_1/n1244 ), .ICI(\mult_x_1/n761 ), .S(
        \mult_x_1/n754 ), .ICO(\mult_x_1/n752 ), .CO(\mult_x_1/n753 ) );
  CMPR42X1TS \mult_x_1/U467  ( .A(\mult_x_1/n751 ), .B(\mult_x_1/n1147 ), .C(
        \mult_x_1/n755 ), .D(\mult_x_1/n1179 ), .ICI(\mult_x_1/n756 ), .S(
        \mult_x_1/n749 ), .ICO(\mult_x_1/n747 ), .CO(\mult_x_1/n748 ) );
  CMPR42X1TS \mult_x_1/U466  ( .A(\mult_x_1/n749 ), .B(\mult_x_1/n752 ), .C(
        \mult_x_1/n1211 ), .D(\mult_x_1/n1243 ), .ICI(\mult_x_1/n753 ), .S(
        \mult_x_1/n746 ), .ICO(\mult_x_1/n744 ), .CO(\mult_x_1/n745 ) );
  CMPR42X1TS \mult_x_1/U464  ( .A(\mult_x_1/n743 ), .B(\mult_x_1/n1146 ), .C(
        \mult_x_1/n747 ), .D(\mult_x_1/n1178 ), .ICI(\mult_x_1/n748 ), .S(
        \mult_x_1/n741 ), .ICO(\mult_x_1/n739 ), .CO(\mult_x_1/n740 ) );
  CMPR42X1TS \mult_x_1/U463  ( .A(\mult_x_1/n741 ), .B(\mult_x_1/n744 ), .C(
        \mult_x_1/n1210 ), .D(\mult_x_1/n1242 ), .ICI(\mult_x_1/n745 ), .S(
        \mult_x_1/n738 ), .ICO(\mult_x_1/n736 ), .CO(\mult_x_1/n737 ) );
  CMPR42X1TS \mult_x_1/U460  ( .A(\mult_x_1/n733 ), .B(\mult_x_1/n739 ), .C(
        \mult_x_1/n1145 ), .D(\mult_x_1/n1177 ), .ICI(\mult_x_1/n740 ), .S(
        \mult_x_1/n731 ), .ICO(\mult_x_1/n729 ), .CO(\mult_x_1/n730 ) );
  CMPR42X1TS \mult_x_1/U459  ( .A(\mult_x_1/n731 ), .B(\mult_x_1/n736 ), .C(
        \mult_x_1/n1209 ), .D(\mult_x_1/n1241 ), .ICI(\mult_x_1/n737 ), .S(
        \mult_x_1/n728 ), .ICO(\mult_x_1/n726 ), .CO(\mult_x_1/n727 ) );
  CMPR42X1TS \mult_x_1/U456  ( .A(\mult_x_1/n723 ), .B(\mult_x_1/n729 ), .C(
        \mult_x_1/n1144 ), .D(\mult_x_1/n1176 ), .ICI(\mult_x_1/n730 ), .S(
        \mult_x_1/n721 ), .ICO(\mult_x_1/n719 ), .CO(\mult_x_1/n720 ) );
  CMPR42X1TS \mult_x_1/U455  ( .A(\mult_x_1/n721 ), .B(\mult_x_1/n726 ), .C(
        \mult_x_1/n1208 ), .D(\mult_x_1/n1240 ), .ICI(\mult_x_1/n727 ), .S(
        \mult_x_1/n718 ), .ICO(\mult_x_1/n716 ), .CO(\mult_x_1/n717 ) );
  CMPR42X1TS \mult_x_1/U452  ( .A(\mult_x_1/n713 ), .B(\mult_x_1/n719 ), .C(
        \mult_x_1/n1143 ), .D(\mult_x_1/n1175 ), .ICI(\mult_x_1/n720 ), .S(
        \mult_x_1/n711 ), .ICO(\mult_x_1/n709 ), .CO(\mult_x_1/n710 ) );
  CMPR42X1TS \mult_x_1/U451  ( .A(\mult_x_1/n711 ), .B(\mult_x_1/n716 ), .C(
        \mult_x_1/n1207 ), .D(\mult_x_1/n1239 ), .ICI(\mult_x_1/n717 ), .S(
        \mult_x_1/n708 ), .ICO(\mult_x_1/n706 ), .CO(\mult_x_1/n707 ) );
  CMPR42X1TS \mult_x_1/U449  ( .A(\mult_x_1/n705 ), .B(\mult_x_1/n1078 ), .C(
        \mult_x_1/n714 ), .D(\mult_x_1/n1110 ), .ICI(\mult_x_1/n712 ), .S(
        \mult_x_1/n703 ), .ICO(\mult_x_1/n701 ), .CO(\mult_x_1/n702 ) );
  CMPR42X1TS \mult_x_1/U448  ( .A(\mult_x_1/n703 ), .B(\mult_x_1/n709 ), .C(
        \mult_x_1/n1142 ), .D(\mult_x_1/n1174 ), .ICI(\mult_x_1/n710 ), .S(
        \mult_x_1/n700 ), .ICO(\mult_x_1/n698 ), .CO(\mult_x_1/n699 ) );
  CMPR42X1TS \mult_x_1/U447  ( .A(\mult_x_1/n700 ), .B(\mult_x_1/n706 ), .C(
        \mult_x_1/n1206 ), .D(\mult_x_1/n1238 ), .ICI(\mult_x_1/n707 ), .S(
        \mult_x_1/n697 ), .ICO(\mult_x_1/n695 ), .CO(\mult_x_1/n696 ) );
  CMPR42X1TS \mult_x_1/U445  ( .A(\mult_x_1/n694 ), .B(\mult_x_1/n1077 ), .C(
        \mult_x_1/n701 ), .D(\mult_x_1/n1109 ), .ICI(\mult_x_1/n702 ), .S(
        \mult_x_1/n692 ), .ICO(\mult_x_1/n690 ), .CO(\mult_x_1/n691 ) );
  CMPR42X1TS \mult_x_1/U444  ( .A(\mult_x_1/n692 ), .B(\mult_x_1/n698 ), .C(
        \mult_x_1/n1141 ), .D(\mult_x_1/n1173 ), .ICI(\mult_x_1/n699 ), .S(
        \mult_x_1/n689 ), .ICO(\mult_x_1/n687 ), .CO(\mult_x_1/n688 ) );
  CMPR42X1TS \mult_x_1/U443  ( .A(\mult_x_1/n689 ), .B(\mult_x_1/n695 ), .C(
        \mult_x_1/n1205 ), .D(\mult_x_1/n1237 ), .ICI(\mult_x_1/n696 ), .S(
        \mult_x_1/n686 ), .ICO(\mult_x_1/n684 ), .CO(\mult_x_1/n685 ) );
  CMPR42X1TS \mult_x_1/U441  ( .A(\mult_x_1/n683 ), .B(\mult_x_1/n1076 ), .C(
        \mult_x_1/n690 ), .D(\mult_x_1/n1108 ), .ICI(\mult_x_1/n691 ), .S(
        \mult_x_1/n681 ), .ICO(\mult_x_1/n679 ), .CO(\mult_x_1/n680 ) );
  CMPR42X1TS \mult_x_1/U440  ( .A(\mult_x_1/n681 ), .B(\mult_x_1/n687 ), .C(
        \mult_x_1/n1140 ), .D(\mult_x_1/n1172 ), .ICI(\mult_x_1/n688 ), .S(
        \mult_x_1/n678 ), .ICO(\mult_x_1/n676 ), .CO(\mult_x_1/n677 ) );
  CMPR42X1TS \mult_x_1/U439  ( .A(\mult_x_1/n678 ), .B(\mult_x_1/n684 ), .C(
        \mult_x_1/n1204 ), .D(\mult_x_1/n1236 ), .ICI(\mult_x_1/n685 ), .S(
        \mult_x_1/n675 ), .ICO(\mult_x_1/n673 ), .CO(\mult_x_1/n674 ) );
  CMPR42X1TS \mult_x_1/U436  ( .A(\mult_x_1/n670 ), .B(\mult_x_1/n679 ), .C(
        \mult_x_1/n1075 ), .D(\mult_x_1/n1107 ), .ICI(\mult_x_1/n680 ), .S(
        \mult_x_1/n668 ), .ICO(\mult_x_1/n666 ), .CO(\mult_x_1/n667 ) );
  CMPR42X1TS \mult_x_1/U435  ( .A(\mult_x_1/n668 ), .B(\mult_x_1/n676 ), .C(
        \mult_x_1/n1139 ), .D(\mult_x_1/n1171 ), .ICI(\mult_x_1/n677 ), .S(
        \mult_x_1/n665 ), .ICO(\mult_x_1/n663 ), .CO(\mult_x_1/n664 ) );
  CMPR42X1TS \mult_x_1/U434  ( .A(\mult_x_1/n665 ), .B(\mult_x_1/n673 ), .C(
        \mult_x_1/n1203 ), .D(\mult_x_1/n1235 ), .ICI(\mult_x_1/n674 ), .S(
        \mult_x_1/n662 ), .ICO(\mult_x_1/n660 ), .CO(\mult_x_1/n661 ) );
  CMPR42X1TS \mult_x_1/U431  ( .A(\mult_x_1/n657 ), .B(\mult_x_1/n666 ), .C(
        \mult_x_1/n1074 ), .D(\mult_x_1/n1106 ), .ICI(\mult_x_1/n667 ), .S(
        \mult_x_1/n655 ), .ICO(\mult_x_1/n653 ), .CO(\mult_x_1/n654 ) );
  CMPR42X1TS \mult_x_1/U430  ( .A(\mult_x_1/n655 ), .B(\mult_x_1/n663 ), .C(
        \mult_x_1/n1138 ), .D(\mult_x_1/n1170 ), .ICI(\mult_x_1/n664 ), .S(
        \mult_x_1/n652 ), .ICO(\mult_x_1/n650 ), .CO(\mult_x_1/n651 ) );
  CMPR42X1TS \mult_x_1/U429  ( .A(\mult_x_1/n652 ), .B(\mult_x_1/n660 ), .C(
        \mult_x_1/n1202 ), .D(\mult_x_1/n1234 ), .ICI(\mult_x_1/n661 ), .S(
        \mult_x_1/n649 ), .ICO(\mult_x_1/n647 ), .CO(\mult_x_1/n648 ) );
  CMPR42X1TS \mult_x_1/U426  ( .A(\mult_x_1/n644 ), .B(\mult_x_1/n653 ), .C(
        \mult_x_1/n1073 ), .D(\mult_x_1/n1105 ), .ICI(\mult_x_1/n654 ), .S(
        \mult_x_1/n642 ), .ICO(\mult_x_1/n640 ), .CO(\mult_x_1/n641 ) );
  CMPR42X1TS \mult_x_1/U425  ( .A(\mult_x_1/n642 ), .B(\mult_x_1/n650 ), .C(
        \mult_x_1/n1137 ), .D(\mult_x_1/n1169 ), .ICI(\mult_x_1/n651 ), .S(
        \mult_x_1/n639 ), .ICO(\mult_x_1/n637 ), .CO(\mult_x_1/n638 ) );
  CMPR42X1TS \mult_x_1/U424  ( .A(\mult_x_1/n639 ), .B(\mult_x_1/n647 ), .C(
        \mult_x_1/n1201 ), .D(\mult_x_1/n1233 ), .ICI(\mult_x_1/n648 ), .S(
        \mult_x_1/n636 ), .ICO(\mult_x_1/n634 ), .CO(\mult_x_1/n635 ) );
  CMPR42X1TS \mult_x_1/U421  ( .A(\mult_x_1/n631 ), .B(\mult_x_1/n640 ), .C(
        \mult_x_1/n1072 ), .D(\mult_x_1/n1104 ), .ICI(\mult_x_1/n641 ), .S(
        \mult_x_1/n628 ), .ICO(\mult_x_1/n626 ), .CO(\mult_x_1/n627 ) );
  CMPR42X1TS \mult_x_1/U420  ( .A(\mult_x_1/n628 ), .B(\mult_x_1/n637 ), .C(
        \mult_x_1/n1136 ), .D(\mult_x_1/n1168 ), .ICI(\mult_x_1/n638 ), .S(
        \mult_x_1/n625 ), .ICO(\mult_x_1/n623 ), .CO(\mult_x_1/n624 ) );
  CMPR42X1TS \mult_x_1/U419  ( .A(\mult_x_1/n625 ), .B(\mult_x_1/n634 ), .C(
        \mult_x_1/n1200 ), .D(\mult_x_1/n1232 ), .ICI(\mult_x_1/n635 ), .S(
        \mult_x_1/n622 ), .ICO(\mult_x_1/n620 ), .CO(\mult_x_1/n621 ) );
  CMPR42X1TS \mult_x_1/U416  ( .A(\mult_x_1/n617 ), .B(\mult_x_1/n626 ), .C(
        \mult_x_1/n1071 ), .D(\mult_x_1/n1103 ), .ICI(\mult_x_1/n627 ), .S(
        \mult_x_1/n614 ), .ICO(\mult_x_1/n612 ), .CO(\mult_x_1/n613 ) );
  CMPR42X1TS \mult_x_1/U415  ( .A(\mult_x_1/n614 ), .B(\mult_x_1/n623 ), .C(
        \mult_x_1/n1135 ), .D(\mult_x_1/n1167 ), .ICI(\mult_x_1/n624 ), .S(
        \mult_x_1/n611 ), .ICO(\mult_x_1/n609 ), .CO(\mult_x_1/n610 ) );
  CMPR42X1TS \mult_x_1/U414  ( .A(\mult_x_1/n611 ), .B(\mult_x_1/n620 ), .C(
        \mult_x_1/n1199 ), .D(\mult_x_1/n1231 ), .ICI(\mult_x_1/n621 ), .S(
        \mult_x_1/n608 ), .ICO(\mult_x_1/n606 ), .CO(\mult_x_1/n607 ) );
  CMPR42X1TS \mult_x_1/U411  ( .A(\mult_x_1/n603 ), .B(\mult_x_1/n612 ), .C(
        \mult_x_1/n1070 ), .D(\mult_x_1/n1102 ), .ICI(\mult_x_1/n613 ), .S(
        \mult_x_1/n600 ), .ICO(\mult_x_1/n598 ), .CO(\mult_x_1/n599 ) );
  CMPR42X1TS \mult_x_1/U410  ( .A(\mult_x_1/n600 ), .B(\mult_x_1/n609 ), .C(
        \mult_x_1/n1134 ), .D(\mult_x_1/n1166 ), .ICI(\mult_x_1/n610 ), .S(
        \mult_x_1/n597 ), .ICO(\mult_x_1/n595 ), .CO(\mult_x_1/n596 ) );
  CMPR42X1TS \mult_x_1/U409  ( .A(\mult_x_1/n597 ), .B(\mult_x_1/n606 ), .C(
        \mult_x_1/n1198 ), .D(n1036), .ICI(\mult_x_1/n607 ), .S(
        \mult_x_1/n594 ), .ICO(\mult_x_1/n592 ), .CO(\mult_x_1/n593 ) );
  CMPR42X1TS \mult_x_1/U406  ( .A(\mult_x_1/n589 ), .B(\mult_x_1/n598 ), .C(
        \mult_x_1/n1069 ), .D(\mult_x_1/n1101 ), .ICI(\mult_x_1/n599 ), .S(
        \mult_x_1/n586 ), .ICO(\mult_x_1/n584 ), .CO(\mult_x_1/n585 ) );
  CMPR42X1TS \mult_x_1/U405  ( .A(\mult_x_1/n586 ), .B(\mult_x_1/n595 ), .C(
        \mult_x_1/n1133 ), .D(\mult_x_1/n1165 ), .ICI(\mult_x_1/n596 ), .S(
        \mult_x_1/n583 ), .ICO(\mult_x_1/n581 ), .CO(\mult_x_1/n582 ) );
  CMPR42X1TS \mult_x_1/U404  ( .A(\mult_x_1/n583 ), .B(\mult_x_1/n592 ), .C(
        \mult_x_1/n1197 ), .D(n1036), .ICI(\mult_x_1/n593 ), .S(
        \mult_x_1/n580 ), .ICO(\mult_x_1/n578 ), .CO(\mult_x_1/n579 ) );
  CMPR42X1TS \mult_x_1/U401  ( .A(\mult_x_1/n575 ), .B(\mult_x_1/n584 ), .C(
        \mult_x_1/n1068 ), .D(\mult_x_1/n1100 ), .ICI(\mult_x_1/n585 ), .S(
        \mult_x_1/n572 ), .ICO(\mult_x_1/n570 ), .CO(\mult_x_1/n571 ) );
  CMPR42X1TS \mult_x_1/U400  ( .A(\mult_x_1/n572 ), .B(\mult_x_1/n581 ), .C(
        \mult_x_1/n1132 ), .D(\mult_x_1/n1164 ), .ICI(\mult_x_1/n582 ), .S(
        \mult_x_1/n569 ), .ICO(\mult_x_1/n567 ), .CO(\mult_x_1/n568 ) );
  CMPR42X1TS \mult_x_1/U399  ( .A(\mult_x_1/n569 ), .B(\mult_x_1/n578 ), .C(
        \mult_x_1/n1196 ), .D(n1036), .ICI(\mult_x_1/n579 ), .S(
        \mult_x_1/n566 ), .ICO(\mult_x_1/n564 ), .CO(\mult_x_1/n565 ) );
  CMPR42X1TS \mult_x_1/U396  ( .A(\mult_x_1/n561 ), .B(\mult_x_1/n570 ), .C(
        \mult_x_1/n1067 ), .D(\mult_x_1/n1099 ), .ICI(\mult_x_1/n571 ), .S(
        \mult_x_1/n558 ), .ICO(\mult_x_1/n556 ), .CO(\mult_x_1/n557 ) );
  CMPR42X1TS \mult_x_1/U395  ( .A(\mult_x_1/n558 ), .B(\mult_x_1/n567 ), .C(
        \mult_x_1/n1131 ), .D(\mult_x_1/n1163 ), .ICI(\mult_x_1/n568 ), .S(
        \mult_x_1/n555 ), .ICO(\mult_x_1/n553 ), .CO(\mult_x_1/n554 ) );
  CMPR42X1TS \mult_x_1/U394  ( .A(\mult_x_1/n555 ), .B(\mult_x_1/n564 ), .C(
        A[8]), .D(n1036), .ICI(\mult_x_1/n565 ), .S(\mult_x_1/n552 ), .ICO(
        \mult_x_1/n550 ), .CO(\mult_x_1/n551 ) );
  CMPR42X1TS \mult_x_1/U391  ( .A(\mult_x_1/n547 ), .B(\mult_x_1/n556 ), .C(
        \mult_x_1/n1066 ), .D(\mult_x_1/n1098 ), .ICI(\mult_x_1/n557 ), .S(
        \mult_x_1/n544 ), .ICO(\mult_x_1/n542 ), .CO(\mult_x_1/n543 ) );
  CMPR42X1TS \mult_x_1/U390  ( .A(\mult_x_1/n544 ), .B(\mult_x_1/n553 ), .C(
        \mult_x_1/n1130 ), .D(\mult_x_1/n1162 ), .ICI(\mult_x_1/n554 ), .S(
        \mult_x_1/n541 ), .ICO(\mult_x_1/n539 ), .CO(\mult_x_1/n540 ) );
  CMPR42X1TS \mult_x_1/U389  ( .A(\mult_x_1/n541 ), .B(\mult_x_1/n550 ), .C(
        A[8]), .D(n1036), .ICI(\mult_x_1/n551 ), .S(\mult_x_1/n538 ), .ICO(
        \mult_x_1/n536 ), .CO(\mult_x_1/n537 ) );
  CMPR42X1TS \mult_x_1/U386  ( .A(\mult_x_1/n546 ), .B(\mult_x_1/n533 ), .C(
        \mult_x_1/n542 ), .D(\mult_x_1/n1065 ), .ICI(\mult_x_1/n1097 ), .S(
        \mult_x_1/n530 ), .ICO(\mult_x_1/n528 ), .CO(\mult_x_1/n529 ) );
  CMPR42X1TS \mult_x_1/U385  ( .A(\mult_x_1/n543 ), .B(\mult_x_1/n530 ), .C(
        \mult_x_1/n539 ), .D(\mult_x_1/n1129 ), .ICI(\mult_x_1/n1161 ), .S(
        \mult_x_1/n527 ), .ICO(\mult_x_1/n525 ), .CO(\mult_x_1/n526 ) );
  CMPR42X1TS \mult_x_1/U384  ( .A(\mult_x_1/n540 ), .B(\mult_x_1/n527 ), .C(
        \mult_x_1/n536 ), .D(A[8]), .ICI(n1036), .S(\mult_x_1/n524 ), .ICO(
        \mult_x_1/n522 ), .CO(\mult_x_1/n523 ) );
  CMPR42X1TS \mult_x_1/U381  ( .A(\mult_x_1/n1032 ), .B(\mult_x_1/n519 ), .C(
        \mult_x_1/n528 ), .D(\mult_x_1/n1064 ), .ICI(\mult_x_1/n529 ), .S(
        \mult_x_1/n516 ), .ICO(\mult_x_1/n514 ), .CO(\mult_x_1/n515 ) );
  CMPR42X1TS \mult_x_1/U380  ( .A(\mult_x_1/n1096 ), .B(\mult_x_1/n516 ), .C(
        \mult_x_1/n525 ), .D(\mult_x_1/n1128 ), .ICI(\mult_x_1/n526 ), .S(
        \mult_x_1/n513 ), .ICO(\mult_x_1/n511 ), .CO(\mult_x_1/n512 ) );
  CMPR42X1TS \mult_x_1/U379  ( .A(A[11]), .B(\mult_x_1/n513 ), .C(
        \mult_x_1/n522 ), .D(A[8]), .ICI(n1036), .S(\mult_x_1/n510 ), .ICO(
        \mult_x_1/n508 ), .CO(\mult_x_1/n509 ) );
  CMPR42X1TS \mult_x_1/U376  ( .A(\mult_x_1/n1031 ), .B(\mult_x_1/n505 ), .C(
        \mult_x_1/n514 ), .D(\mult_x_1/n1063 ), .ICI(\mult_x_1/n515 ), .S(
        \mult_x_1/n502 ), .ICO(\mult_x_1/n500 ), .CO(\mult_x_1/n501 ) );
  CMPR42X1TS \mult_x_1/U375  ( .A(\mult_x_1/n1095 ), .B(\mult_x_1/n502 ), .C(
        \mult_x_1/n511 ), .D(\mult_x_1/n1127 ), .ICI(\mult_x_1/n512 ), .S(
        \mult_x_1/n499 ), .ICO(\mult_x_1/n497 ), .CO(\mult_x_1/n498 ) );
  CMPR42X1TS \mult_x_1/U374  ( .A(A[11]), .B(\mult_x_1/n499 ), .C(
        \mult_x_1/n508 ), .D(A[8]), .ICI(n1036), .S(\mult_x_1/n496 ), .ICO(
        \mult_x_1/n494 ), .CO(\mult_x_1/n495 ) );
  CMPR42X1TS \mult_x_1/U371  ( .A(\mult_x_1/n491 ), .B(n1034), .C(
        \mult_x_1/n1030 ), .D(\mult_x_1/n500 ), .ICI(\mult_x_1/n1062 ), .S(
        \mult_x_1/n488 ), .ICO(\mult_x_1/n486 ), .CO(\mult_x_1/n487 ) );
  CMPR42X1TS \mult_x_1/U370  ( .A(\mult_x_1/n488 ), .B(\mult_x_1/n501 ), .C(
        \mult_x_1/n1094 ), .D(\mult_x_1/n497 ), .ICI(\mult_x_1/n1126 ), .S(
        \mult_x_1/n485 ), .ICO(\mult_x_1/n483 ), .CO(\mult_x_1/n484 ) );
  CMPR42X1TS \mult_x_1/U369  ( .A(\mult_x_1/n485 ), .B(\mult_x_1/n498 ), .C(
        A[11]), .D(\mult_x_1/n494 ), .ICI(A[8]), .S(\mult_x_1/n482 ), .ICO(
        \mult_x_1/n480 ), .CO(\mult_x_1/n481 ) );
  CMPR42X1TS \mult_x_1/U366  ( .A(B[14]), .B(\mult_x_1/n464 ), .C(
        \mult_x_1/n486 ), .D(\mult_x_1/n1029 ), .ICI(\mult_x_1/n487 ), .S(
        \mult_x_1/n475 ), .ICO(\mult_x_1/n473 ), .CO(\mult_x_1/n474 ) );
  CMPR42X1TS \mult_x_1/U365  ( .A(\mult_x_1/n1061 ), .B(\mult_x_1/n475 ), .C(
        \mult_x_1/n483 ), .D(\mult_x_1/n1093 ), .ICI(\mult_x_1/n484 ), .S(
        \mult_x_1/n472 ), .ICO(\mult_x_1/n470 ), .CO(\mult_x_1/n471 ) );
  CMPR42X1TS \mult_x_1/U364  ( .A(A[14]), .B(\mult_x_1/n472 ), .C(
        \mult_x_1/n480 ), .D(A[11]), .ICI(A[8]), .S(\mult_x_1/n469 ), .ICO(
        \mult_x_1/n467 ), .CO(\mult_x_1/n468 ) );
  CMPR42X1TS \mult_x_1/U361  ( .A(B[15]), .B(\mult_x_1/n464 ), .C(
        \mult_x_1/n473 ), .D(\mult_x_1/n1028 ), .ICI(\mult_x_1/n474 ), .S(
        \mult_x_1/n461 ), .ICO(\mult_x_1/n459 ), .CO(\mult_x_1/n460 ) );
  CMPR42X1TS \mult_x_1/U360  ( .A(\mult_x_1/n1060 ), .B(\mult_x_1/n461 ), .C(
        \mult_x_1/n470 ), .D(\mult_x_1/n1092 ), .ICI(\mult_x_1/n471 ), .S(
        \mult_x_1/n458 ), .ICO(\mult_x_1/n456 ), .CO(\mult_x_1/n457 ) );
  CMPR42X1TS \mult_x_1/U359  ( .A(A[14]), .B(\mult_x_1/n458 ), .C(
        \mult_x_1/n467 ), .D(A[11]), .ICI(A[8]), .S(\mult_x_1/n455 ), .ICO(
        \mult_x_1/n453 ), .CO(\mult_x_1/n454 ) );
  CMPR42X1TS \mult_x_1/U357  ( .A(\mult_x_1/n452 ), .B(\mult_x_1/n463 ), .C(
        B[16]), .D(\mult_x_1/n459 ), .ICI(\mult_x_1/n1027 ), .S(
        \mult_x_1/n450 ), .ICO(\mult_x_1/n448 ), .CO(\mult_x_1/n449 ) );
  CMPR42X1TS \mult_x_1/U356  ( .A(\mult_x_1/n450 ), .B(\mult_x_1/n460 ), .C(
        \mult_x_1/n1059 ), .D(\mult_x_1/n456 ), .ICI(\mult_x_1/n1091 ), .S(
        \mult_x_1/n447 ), .ICO(\mult_x_1/n445 ), .CO(\mult_x_1/n446 ) );
  CMPR42X1TS \mult_x_1/U355  ( .A(\mult_x_1/n447 ), .B(\mult_x_1/n457 ), .C(
        A[14]), .D(\mult_x_1/n453 ), .ICI(A[11]), .S(\mult_x_1/n444 ), .ICO(
        \mult_x_1/n442 ), .CO(\mult_x_1/n443 ) );
  CMPR42X1TS \mult_x_1/U351  ( .A(\mult_x_1/n449 ), .B(\mult_x_1/n438 ), .C(
        \mult_x_1/n445 ), .D(\mult_x_1/n1058 ), .ICI(A[17]), .S(
        \mult_x_1/n435 ), .ICO(\mult_x_1/n433 ), .CO(\mult_x_1/n434 ) );
  CMPR42X1TS \mult_x_1/U350  ( .A(\mult_x_1/n446 ), .B(\mult_x_1/n435 ), .C(
        \mult_x_1/n442 ), .D(A[14]), .ICI(A[11]), .S(\mult_x_1/n432 ), .ICO(
        \mult_x_1/n430 ), .CO(\mult_x_1/n431 ) );
  CMPR42X1TS \mult_x_1/U346  ( .A(\mult_x_1/n1025 ), .B(\mult_x_1/n425 ), .C(
        \mult_x_1/n433 ), .D(\mult_x_1/n1057 ), .ICI(\mult_x_1/n434 ), .S(
        \mult_x_1/n422 ), .ICO(\mult_x_1/n420 ), .CO(\mult_x_1/n421 ) );
  CMPR42X1TS \mult_x_1/U345  ( .A(A[17]), .B(\mult_x_1/n422 ), .C(
        \mult_x_1/n430 ), .D(A[14]), .ICI(A[11]), .S(\mult_x_1/n419 ), .ICO(
        \mult_x_1/n417 ), .CO(\mult_x_1/n418 ) );
  CMPR42X1TS \mult_x_1/U342  ( .A(\mult_x_1/n414 ), .B(\mult_x_1/n424 ), .C(
        \mult_x_1/n1024 ), .D(\mult_x_1/n420 ), .ICI(\mult_x_1/n1056 ), .S(
        \mult_x_1/n411 ), .ICO(\mult_x_1/n409 ), .CO(\mult_x_1/n410 ) );
  CMPR42X1TS \mult_x_1/U341  ( .A(\mult_x_1/n411 ), .B(\mult_x_1/n421 ), .C(
        A[17]), .D(\mult_x_1/n417 ), .ICI(A[14]), .S(\mult_x_1/n408 ), .ICO(
        \mult_x_1/n406 ), .CO(\mult_x_1/n407 ) );
  CMPR42X1TS \mult_x_1/U338  ( .A(\mult_x_1/n413 ), .B(\mult_x_1/n404 ), .C(
        \mult_x_1/n409 ), .D(\mult_x_1/n1023 ), .ICI(A[20]), .S(
        \mult_x_1/n401 ), .ICO(\mult_x_1/n399 ), .CO(\mult_x_1/n400 ) );
  CMPR42X1TS \mult_x_1/U337  ( .A(\mult_x_1/n410 ), .B(\mult_x_1/n401 ), .C(
        \mult_x_1/n406 ), .D(A[17]), .ICI(A[14]), .S(\mult_x_1/n398 ), .ICO(
        \mult_x_1/n396 ), .CO(\mult_x_1/n397 ) );
  CMPR42X1TS \mult_x_1/U334  ( .A(B[21]), .B(\mult_x_1/n404 ), .C(
        \mult_x_1/n399 ), .D(\mult_x_1/n1022 ), .ICI(\mult_x_1/n400 ), .S(
        \mult_x_1/n390 ), .ICO(\mult_x_1/n388 ), .CO(\mult_x_1/n389 ) );
  CMPR42X1TS \mult_x_1/U333  ( .A(A[20]), .B(\mult_x_1/n390 ), .C(
        \mult_x_1/n396 ), .D(A[17]), .ICI(A[14]), .S(\mult_x_1/n387 ), .ICO(
        \mult_x_1/n385 ), .CO(\mult_x_1/n386 ) );
  CMPR42X1TS \mult_x_1/U331  ( .A(n1035), .B(B[20]), .C(B[22]), .D(
        \mult_x_1/n388 ), .ICI(\mult_x_1/n1021 ), .S(\mult_x_1/n382 ), .ICO(
        \mult_x_1/n363 ), .CO(\mult_x_1/n381 ) );
  CMPR42X1TS \mult_x_1/U330  ( .A(\mult_x_1/n382 ), .B(\mult_x_1/n389 ), .C(
        A[20]), .D(\mult_x_1/n385 ), .ICI(A[17]), .S(\mult_x_1/n379 ), .ICO(
        \mult_x_1/n377 ), .CO(\mult_x_1/n378 ) );
  CMPR42X1TS \mult_x_1/U326  ( .A(\mult_x_1/n381 ), .B(\mult_x_1/n373 ), .C(
        \mult_x_1/n377 ), .D(A[20]), .ICI(A[17]), .S(\mult_x_1/n370 ), .ICO(
        \mult_x_1/n368 ), .CO(\mult_x_1/n369 ) );
  NAND3X2TS U1 ( .A(n523), .B(n492), .C(n524), .Y(n1017) );
  OR3X2TS U2 ( .A(n96), .B(n135), .C(n95), .Y(n93) );
  NAND3X2TS U3 ( .A(n354), .B(n163), .C(n355), .Y(n1011) );
  NAND2X2TS U4 ( .A(n403), .B(n451), .Y(n404) );
  NAND2X2TS U5 ( .A(n663), .B(n651), .Y(n652) );
  NAND2X2TS U6 ( .A(n87), .B(n81), .Y(n80) );
  CLKAND2X2TS U7 ( .A(A[0]), .B(n11), .Y(n5) );
  INVX2TS U8 ( .A(A[20]), .Y(n917) );
  ADDFX1TS U9 ( .A(n819), .B(n376), .CI(n375), .CO(n372), .S(n377) );
  ADDFX1TS U10 ( .A(n885), .B(n385), .CI(n384), .CO(n387), .S(n386) );
  ADDFX1TS U11 ( .A(n864), .B(n391), .CI(n390), .CO(n369), .S(n392) );
  ADDFX1TS U12 ( .A(n817), .B(n394), .CI(n393), .CO(n375), .S(n395) );
  ADDFX1TS U13 ( .A(n882), .B(n379), .CI(n378), .CO(n381), .S(n380) );
  ADDFX1TS U14 ( .A(n884), .B(n382), .CI(n381), .CO(n384), .S(n383) );
  ADDFX1TS U15 ( .A(n921), .B(B[10]), .CI(A[2]), .CO(n319), .S(\mult_x_1/n533 ) );
  ADDFX1TS U16 ( .A(A[2]), .B(B[11]), .CI(n319), .CO(n314), .S(\mult_x_1/n519 ) );
  ADDFX1TS U17 ( .A(A[2]), .B(B[12]), .CI(n314), .CO(n1034), .S(
        \mult_x_1/n505 ) );
  ADDFX1TS U18 ( .A(n821), .B(n373), .CI(n372), .CO(n378), .S(n374) );
  ADDFX1TS U19 ( .A(n852), .B(n388), .CI(n387), .CO(n390), .S(n389) );
  ADDFX1TS U20 ( .A(n877), .B(n370), .CI(n369), .CO(n353), .S(n371) );
  ADDFX1TS U21 ( .A(n905), .B(n298), .CI(n297), .CO(n300), .S(n299) );
  ADDFX1TS U22 ( .A(n988), .B(n301), .CI(n300), .CO(n290), .S(n302) );
  ADDFX1TS U23 ( .A(n992), .B(A[11]), .CI(n283), .CO(n212), .S(n221) );
  ADDFX1TS U24 ( .A(B[7]), .B(B[8]), .CI(n72), .CO(n68), .S(n332) );
  ADDFX1TS U25 ( .A(B[17]), .B(B[18]), .CI(n30), .CO(n26), .S(n990) );
  ADDFX1TS U26 ( .A(B[4]), .B(B[5]), .CI(n111), .CO(n125), .S(n341) );
  ADDFX1TS U27 ( .A(B[5]), .B(B[6]), .CI(n125), .CO(n118), .S(n338) );
  ADDFX1TS U28 ( .A(B[6]), .B(B[7]), .CI(n118), .CO(n72), .S(n335) );
  ADDFX1TS U29 ( .A(B[9]), .B(B[10]), .CI(n64), .CO(n60), .S(n326) );
  ADDFX1TS U30 ( .A(B[10]), .B(B[11]), .CI(n60), .CO(n56), .S(n323) );
  ADDFX1TS U31 ( .A(B[11]), .B(B[12]), .CI(n56), .CO(n52), .S(n320) );
  ADDFX1TS U32 ( .A(B[12]), .B(B[13]), .CI(n52), .CO(n48), .S(n313) );
  ADDFX1TS U33 ( .A(B[13]), .B(B[14]), .CI(n48), .CO(n44), .S(n975) );
  ADDFX1TS U34 ( .A(B[14]), .B(B[15]), .CI(n44), .CO(n39), .S(n979) );
  ADDFX1TS U35 ( .A(B[15]), .B(B[16]), .CI(n39), .CO(n34), .S(n40) );
  ADDFX1TS U36 ( .A(B[16]), .B(B[17]), .CI(n34), .CO(n30), .S(n35) );
  ADDFX1TS U37 ( .A(B[18]), .B(B[19]), .CI(n26), .CO(n22), .S(n994) );
  ADDFX1TS U38 ( .A(n560), .B(n559), .CI(n558), .CO(n575), .S(n516) );
  ADDFX1TS U39 ( .A(B[19]), .B(B[20]), .CI(n22), .CO(n18), .S(n287) );
  ADDFX1TS U40 ( .A(n576), .B(n575), .CI(n574), .CO(n564), .S(n577) );
  ADDFX1TS U41 ( .A(B[21]), .B(B[20]), .CI(n18), .CO(n14), .S(n998) );
  ADDFX1TS U42 ( .A(B[3]), .B(B[4]), .CI(n94), .CO(n111), .S(n350) );
  ADDFX1TS U43 ( .A(B[8]), .B(B[9]), .CI(n68), .CO(n64), .S(n329) );
  ADDFX1TS U44 ( .A(B[21]), .B(B[22]), .CI(n14), .CO(n10), .S(n1004) );
  ADDFX1TS U45 ( .A(B[2]), .B(B[3]), .CI(n105), .CO(n94), .S(n349) );
  ADDFX1TS U46 ( .A(n689), .B(n688), .CI(n687), .CO(n749), .S(n682) );
  ADDFX1TS U47 ( .A(n750), .B(n749), .CI(n748), .CO(n693), .S(n751) );
  ADDFX1TS U48 ( .A(n912), .B(n911), .CI(n910), .CO(n913), .S(n185) );
  ADDFX1TS U49 ( .A(n117), .B(n116), .CI(n115), .CO(n911), .S(n182) );
  ADDFX1TS U50 ( .A(n260), .B(n1027), .CI(n259), .CO(n262), .S(n261) );
  ADDFX1TS U51 ( .A(n272), .B(n1027), .CI(n271), .CO(n274), .S(n273) );
  ADDFX1TS U52 ( .A(n278), .B(n1027), .CI(n277), .CO(n280), .S(n279) );
  ADDFX1TS U53 ( .A(n317), .B(n316), .CI(n315), .CO(n362), .S(n318) );
  ADDFX1TS U54 ( .A(n487), .B(n486), .CI(n485), .CO(n505), .S(n488) );
  ADDFX1TS U55 ( .A(n649), .B(n648), .CI(n647), .CO(n659), .S(n650) );
  ADDFX1TS U56 ( .A(n249), .B(n248), .CI(n247), .CO(n251), .S(n250) );
  ADDFX1TS U57 ( .A(n257), .B(n256), .CI(n255), .CO(n259), .S(n258) );
  ADDFX1TS U58 ( .A(n266), .B(n1027), .CI(n265), .CO(n268), .S(n267) );
  ADDFX1TS U59 ( .A(n269), .B(n1027), .CI(n268), .CO(n271), .S(n270) );
  ADDFX1TS U60 ( .A(n293), .B(n292), .CI(n291), .CO(n303), .S(n294) );
  ADDFX1TS U61 ( .A(n305), .B(n304), .CI(n303), .CO(n307), .S(n306) );
  ADDFX1TS U62 ( .A(n309), .B(n308), .CI(n307), .CO(n315), .S(n310) );
  ADDFX1TS U63 ( .A(n364), .B(n363), .CI(n362), .CO(n399), .S(n365) );
  ADDFX1TS U64 ( .A(n419), .B(n418), .CI(n417), .CO(n461), .S(n420) );
  ADDFX1TS U65 ( .A(n463), .B(n462), .CI(n461), .CO(n485), .S(n464) );
  ADDFX1TS U66 ( .A(n507), .B(n506), .CI(n505), .CO(n632), .S(n508) );
  ADDFX1TS U67 ( .A(n253), .B(n252), .CI(n251), .CO(n255), .S(n254) );
  ADDFX1TS U68 ( .A(n263), .B(n1027), .CI(n262), .CO(n265), .S(n264) );
  ADDFX1TS U69 ( .A(n275), .B(n1027), .CI(n274), .CO(n277), .S(n276) );
  ADDFX1TS U70 ( .A(n1027), .B(n281), .CI(n280), .CO(n291), .S(n282) );
  ADDFX1TS U71 ( .A(n401), .B(n400), .CI(n399), .CO(n417), .S(n402) );
  ADDFX1TS U72 ( .A(n634), .B(n633), .CI(n632), .CO(n647), .S(n635) );
  ADDFX1TS U73 ( .A(n805), .B(n804), .CI(n803), .CO(n825), .S(n806) );
  ADDFX1TS U74 ( .A(n186), .B(n185), .CI(n184), .CO(n188), .S(n187) );
  ADDFX1TS U75 ( .A(n228), .B(n227), .CI(n226), .CO(n230), .S(n229) );
  ADDFX1TS U76 ( .A(n174), .B(n173), .CI(n172), .CO(n176), .S(n175) );
  ADDFX1TS U77 ( .A(n178), .B(n177), .CI(n176), .CO(n180), .S(n179) );
  ADDFX1TS U78 ( .A(n182), .B(n181), .CI(n180), .CO(n184), .S(n183) );
  ADDFX1TS U79 ( .A(n194), .B(n193), .CI(n192), .CO(n196), .S(n195) );
  ADDFX1TS U80 ( .A(n198), .B(n197), .CI(n196), .CO(n200), .S(n199) );
  ADDFX1TS U81 ( .A(n202), .B(n201), .CI(n200), .CO(n204), .S(n203) );
  ADDFX1TS U82 ( .A(n206), .B(n205), .CI(n204), .CO(n208), .S(n207) );
  ADDFX1TS U83 ( .A(n210), .B(n209), .CI(n208), .CO(n213), .S(n211) );
  ADDFX1TS U84 ( .A(n215), .B(n214), .CI(n213), .CO(n217), .S(n216) );
  ADDFX1TS U85 ( .A(n219), .B(n218), .CI(n217), .CO(n222), .S(n220) );
  ADDFX1TS U86 ( .A(n224), .B(n223), .CI(n222), .CO(n226), .S(n225) );
  ADDFX1TS U87 ( .A(n232), .B(n231), .CI(n230), .CO(n234), .S(n233) );
  ADDFX1TS U88 ( .A(n236), .B(n235), .CI(n234), .CO(n238), .S(n237) );
  ADDFX1TS U89 ( .A(n240), .B(n239), .CI(n238), .CO(n243), .S(n241) );
  ADDFX1TS U90 ( .A(n245), .B(n244), .CI(n243), .CO(n247), .S(n246) );
  ADDFX1TS U91 ( .A(n170), .B(n922), .CI(n169), .CO(n172), .S(n171) );
  ADDFX1TS U92 ( .A(n190), .B(n189), .CI(n188), .CO(n192), .S(n191) );
  ADDFX1TS U93 ( .A(n661), .B(n660), .CI(n659), .CO(n803), .S(n662) );
  ADDFX1TS U94 ( .A(A[17]), .B(A[20]), .CI(n159), .CO(n918), .S(n4) );
  ADDFX1TS U95 ( .A(n827), .B(n826), .CI(n825), .CO(n158), .S(n828) );
  ADDFX1TS U96 ( .A(n917), .B(n3), .CI(A[17]), .CO(n1), .S(n2) );
  ADDFX1TS U97 ( .A(n917), .B(n916), .CI(n915), .CO(n914), .S(Product[50]) );
  ADDFX1TS U98 ( .A(n920), .B(n919), .CI(n918), .CO(n915), .S(Product[49]) );
  NOR2XLTS U99 ( .A(\mult_x_1/n363 ), .B(\mult_x_1/n368 ), .Y(n3) );
  INVX2TS U100 ( .A(n1), .Y(n916) );
  INVX2TS U101 ( .A(n2), .Y(n920) );
  INVX2TS U102 ( .A(\mult_x_1/n369 ), .Y(n827) );
  AO21XLTS U103 ( .A0(\mult_x_1/n368 ), .A1(\mult_x_1/n363 ), .B0(n3), .Y(n159) );
  INVX2TS U104 ( .A(n4), .Y(n826) );
  INVX2TS U105 ( .A(\mult_x_1/n378 ), .Y(n805) );
  INVX2TS U106 ( .A(\mult_x_1/n370 ), .Y(n804) );
  INVX2TS U107 ( .A(\mult_x_1/n386 ), .Y(n661) );
  INVX2TS U108 ( .A(\mult_x_1/n379 ), .Y(n660) );
  INVX2TS U109 ( .A(\mult_x_1/n397 ), .Y(n649) );
  INVX2TS U110 ( .A(\mult_x_1/n387 ), .Y(n648) );
  INVX2TS U111 ( .A(\mult_x_1/n407 ), .Y(n634) );
  INVX2TS U112 ( .A(\mult_x_1/n398 ), .Y(n633) );
  INVX2TS U113 ( .A(\mult_x_1/n418 ), .Y(n507) );
  INVX2TS U114 ( .A(\mult_x_1/n408 ), .Y(n506) );
  INVX2TS U115 ( .A(\mult_x_1/n431 ), .Y(n487) );
  INVX2TS U116 ( .A(\mult_x_1/n419 ), .Y(n486) );
  INVX2TS U117 ( .A(\mult_x_1/n443 ), .Y(n463) );
  INVX2TS U118 ( .A(\mult_x_1/n432 ), .Y(n462) );
  INVX2TS U119 ( .A(\mult_x_1/n454 ), .Y(n419) );
  INVX2TS U120 ( .A(\mult_x_1/n444 ), .Y(n418) );
  INVX2TS U121 ( .A(\mult_x_1/n468 ), .Y(n401) );
  INVX2TS U122 ( .A(\mult_x_1/n455 ), .Y(n400) );
  INVX2TS U123 ( .A(\mult_x_1/n481 ), .Y(n364) );
  INVX2TS U124 ( .A(\mult_x_1/n469 ), .Y(n363) );
  INVX2TS U125 ( .A(\mult_x_1/n495 ), .Y(n317) );
  INVX2TS U126 ( .A(\mult_x_1/n482 ), .Y(n316) );
  INVX2TS U127 ( .A(\mult_x_1/n509 ), .Y(n309) );
  INVX2TS U128 ( .A(\mult_x_1/n496 ), .Y(n308) );
  INVX2TS U129 ( .A(\mult_x_1/n523 ), .Y(n305) );
  INVX2TS U130 ( .A(\mult_x_1/n510 ), .Y(n304) );
  INVX2TS U131 ( .A(\mult_x_1/n537 ), .Y(n293) );
  INVX2TS U132 ( .A(\mult_x_1/n524 ), .Y(n292) );
  INVX2TS U133 ( .A(A[2]), .Y(n1027) );
  INVX2TS U134 ( .A(\mult_x_1/n538 ), .Y(n281) );
  INVX2TS U135 ( .A(\mult_x_1/n552 ), .Y(n278) );
  INVX2TS U136 ( .A(\mult_x_1/n566 ), .Y(n275) );
  INVX2TS U137 ( .A(\mult_x_1/n580 ), .Y(n272) );
  INVX2TS U138 ( .A(\mult_x_1/n594 ), .Y(n269) );
  INVX2TS U139 ( .A(\mult_x_1/n608 ), .Y(n266) );
  INVX2TS U140 ( .A(\mult_x_1/n622 ), .Y(n263) );
  INVX2TS U141 ( .A(\mult_x_1/n636 ), .Y(n260) );
  INVX2TS U142 ( .A(\mult_x_1/n649 ), .Y(n257) );
  AOI2BB2XLTS U143 ( .B0(A[2]), .B1(A[1]), .A0N(A[1]), .A1N(A[2]), .Y(n11) );
  INVX2TS U144 ( .A(B[2]), .Y(n819) );
  INVX2TS U145 ( .A(B[0]), .Y(n928) );
  INVX2TS U146 ( .A(B[1]), .Y(n817) );
  AOI21X1TS U147 ( .A0(n819), .A1(n928), .B0(n817), .Y(n105) );
  NOR2X1TS U148 ( .A(B[22]), .B(n10), .Y(n1022) );
  INVX2TS U149 ( .A(n1022), .Y(n1009) );
  NAND2X1TS U150 ( .A(n5), .B(n1009), .Y(n7) );
  NOR3XLTS U151 ( .A(A[0]), .B(A[1]), .C(n1027), .Y(n146) );
  INVX2TS U152 ( .A(n146), .Y(n152) );
  INVX2TS U153 ( .A(n7), .Y(n6) );
  AOI32X1TS U154 ( .A0(A[2]), .A1(n7), .A2(n152), .B0(n1027), .B1(n6), .Y(n256) );
  INVX2TS U155 ( .A(\mult_x_1/n662 ), .Y(n253) );
  INVX2TS U156 ( .A(A[0]), .Y(n142) );
  NAND2X2TS U157 ( .A(A[1]), .B(n142), .Y(n154) );
  INVX2TS U158 ( .A(n154), .Y(n143) );
  INVX2TS U159 ( .A(B[22]), .Y(n1001) );
  INVX2TS U160 ( .A(n5), .Y(n151) );
  OAI22X1TS U161 ( .A0(n152), .A1(n1001), .B0(n151), .B1(n1009), .Y(n9) );
  OAI21XLTS U162 ( .A0(n143), .A1(n9), .B0(A[2]), .Y(n8) );
  OAI31X1TS U163 ( .A0(n143), .A1(A[2]), .A2(n9), .B0(n8), .Y(n252) );
  INVX2TS U164 ( .A(\mult_x_1/n675 ), .Y(n249) );
  AOI21X1TS U165 ( .A0(n10), .A1(B[22]), .B0(n1022), .Y(n967) );
  AOI22X1TS U166 ( .A0(n143), .A1(B[22]), .B0(n146), .B1(B[21]), .Y(n12) );
  NOR2XLTS U167 ( .A(n142), .B(n11), .Y(n144) );
  INVX2TS U168 ( .A(n144), .Y(n153) );
  OAI211XLTS U169 ( .A0(n967), .A1(n151), .B0(n12), .C0(n153), .Y(n13) );
  XNOR2X1TS U170 ( .A(A[2]), .B(n13), .Y(n248) );
  INVX2TS U171 ( .A(\mult_x_1/n686 ), .Y(n245) );
  INVX2TS U172 ( .A(B[20]), .Y(\mult_x_1/n404 ) );
  INVX2TS U173 ( .A(n1004), .Y(n835) );
  OAI22X1TS U174 ( .A0(n152), .A1(\mult_x_1/n404 ), .B0(n151), .B1(n835), .Y(
        n17) );
  INVX2TS U175 ( .A(B[21]), .Y(n996) );
  OAI22X1TS U176 ( .A0(n153), .A1(n1001), .B0(n154), .B1(n996), .Y(n16) );
  OAI21XLTS U177 ( .A0(n17), .A1(n16), .B0(A[2]), .Y(n15) );
  OAI31X1TS U178 ( .A0(n17), .A1(A[2]), .A2(n16), .B0(n15), .Y(n244) );
  INVX2TS U179 ( .A(\mult_x_1/n697 ), .Y(n240) );
  INVX2TS U180 ( .A(B[19]), .Y(n992) );
  INVX2TS U181 ( .A(n998), .Y(n831) );
  OAI22X1TS U182 ( .A0(n152), .A1(n992), .B0(n151), .B1(n831), .Y(n21) );
  OAI22X1TS U183 ( .A0(n153), .A1(n996), .B0(n154), .B1(\mult_x_1/n404 ), .Y(
        n20) );
  OAI21XLTS U184 ( .A0(n21), .A1(n20), .B0(A[2]), .Y(n19) );
  OAI31X1TS U185 ( .A0(n21), .A1(A[2]), .A2(n20), .B0(n19), .Y(n239) );
  INVX2TS U186 ( .A(\mult_x_1/n708 ), .Y(n236) );
  INVX2TS U187 ( .A(B[18]), .Y(n988) );
  INVX2TS U188 ( .A(n287), .Y(n889) );
  OAI22X1TS U189 ( .A0(n152), .A1(n988), .B0(n151), .B1(n889), .Y(n25) );
  OAI22X1TS U190 ( .A0(n153), .A1(\mult_x_1/n404 ), .B0(n154), .B1(n992), .Y(
        n24) );
  OAI21XLTS U191 ( .A0(n25), .A1(n24), .B0(A[2]), .Y(n23) );
  OAI31X1TS U192 ( .A0(n25), .A1(A[2]), .A2(n24), .B0(n23), .Y(n235) );
  INVX2TS U193 ( .A(\mult_x_1/n718 ), .Y(n232) );
  INVX2TS U194 ( .A(B[17]), .Y(n905) );
  INVX2TS U195 ( .A(n994), .Y(n856) );
  OAI22X1TS U196 ( .A0(n152), .A1(n905), .B0(n151), .B1(n856), .Y(n29) );
  OAI22X1TS U197 ( .A0(n153), .A1(n992), .B0(n154), .B1(n988), .Y(n28) );
  OAI21XLTS U198 ( .A0(n29), .A1(n28), .B0(A[2]), .Y(n27) );
  OAI31X1TS U199 ( .A0(n29), .A1(A[2]), .A2(n28), .B0(n27), .Y(n231) );
  INVX2TS U200 ( .A(\mult_x_1/n728 ), .Y(n228) );
  INVX2TS U201 ( .A(B[16]), .Y(n903) );
  INVX2TS U202 ( .A(n990), .Y(n869) );
  OAI22X1TS U203 ( .A0(n152), .A1(n903), .B0(n151), .B1(n869), .Y(n33) );
  OAI22X1TS U204 ( .A0(n153), .A1(n988), .B0(n154), .B1(n905), .Y(n32) );
  OAI21XLTS U205 ( .A0(n33), .A1(n32), .B0(A[2]), .Y(n31) );
  OAI31X1TS U206 ( .A0(n33), .A1(A[2]), .A2(n32), .B0(n31), .Y(n227) );
  INVX2TS U207 ( .A(\mult_x_1/n738 ), .Y(n224) );
  INVX2TS U208 ( .A(B[15]), .Y(n977) );
  INVX2TS U209 ( .A(n35), .Y(n985) );
  OAI22X1TS U210 ( .A0(n152), .A1(n977), .B0(n151), .B1(n985), .Y(n38) );
  OAI22X1TS U211 ( .A0(n153), .A1(n905), .B0(n154), .B1(n903), .Y(n37) );
  OAI21XLTS U212 ( .A0(n38), .A1(n37), .B0(A[2]), .Y(n36) );
  OAI31X1TS U213 ( .A0(n38), .A1(A[2]), .A2(n37), .B0(n36), .Y(n223) );
  INVX2TS U214 ( .A(\mult_x_1/n746 ), .Y(n219) );
  INVX2TS U215 ( .A(B[14]), .Y(n973) );
  INVX2TS U216 ( .A(n40), .Y(n981) );
  OAI22X1TS U217 ( .A0(n152), .A1(n973), .B0(n151), .B1(n981), .Y(n43) );
  OAI22X1TS U218 ( .A0(n153), .A1(n903), .B0(n154), .B1(n977), .Y(n42) );
  OAI21XLTS U219 ( .A0(n43), .A1(n42), .B0(A[2]), .Y(n41) );
  OAI31X1TS U220 ( .A0(n43), .A1(A[2]), .A2(n42), .B0(n41), .Y(n218) );
  INVX2TS U221 ( .A(\mult_x_1/n754 ), .Y(n215) );
  INVX2TS U222 ( .A(B[13]), .Y(n1030) );
  INVX2TS U223 ( .A(n979), .Y(n860) );
  OAI22X1TS U224 ( .A0(n152), .A1(n1030), .B0(n151), .B1(n860), .Y(n47) );
  OAI22X1TS U225 ( .A0(n153), .A1(n977), .B0(n154), .B1(n973), .Y(n46) );
  OAI21XLTS U226 ( .A0(n47), .A1(n46), .B0(A[2]), .Y(n45) );
  OAI31X1TS U227 ( .A0(n47), .A1(A[2]), .A2(n46), .B0(n45), .Y(n214) );
  INVX2TS U228 ( .A(\mult_x_1/n762 ), .Y(n210) );
  INVX2TS U229 ( .A(B[12]), .Y(n896) );
  INVX2TS U230 ( .A(n975), .Y(n873) );
  OAI22X1TS U231 ( .A0(n152), .A1(n896), .B0(n151), .B1(n873), .Y(n51) );
  OAI22X1TS U232 ( .A0(n153), .A1(n973), .B0(n154), .B1(n1030), .Y(n50) );
  OAI21XLTS U233 ( .A0(n51), .A1(n50), .B0(A[2]), .Y(n49) );
  OAI31X1TS U234 ( .A0(n51), .A1(A[2]), .A2(n50), .B0(n49), .Y(n209) );
  INVX2TS U235 ( .A(\mult_x_1/n769 ), .Y(n206) );
  INVX2TS U236 ( .A(B[11]), .Y(n895) );
  INVX2TS U237 ( .A(n313), .Y(n839) );
  OAI22X1TS U238 ( .A0(n152), .A1(n895), .B0(n151), .B1(n839), .Y(n55) );
  OAI22X1TS U239 ( .A0(n153), .A1(n1030), .B0(n154), .B1(n896), .Y(n54) );
  OAI21XLTS U240 ( .A0(n55), .A1(n54), .B0(A[2]), .Y(n53) );
  OAI31X1TS U241 ( .A0(n55), .A1(A[2]), .A2(n54), .B0(n53), .Y(n205) );
  INVX2TS U242 ( .A(\mult_x_1/n776 ), .Y(n202) );
  INVX2TS U243 ( .A(B[10]), .Y(n893) );
  INVX2TS U244 ( .A(n320), .Y(n894) );
  OAI22X1TS U245 ( .A0(n152), .A1(n893), .B0(n151), .B1(n894), .Y(n59) );
  OAI22X1TS U246 ( .A0(n153), .A1(n896), .B0(n154), .B1(n895), .Y(n58) );
  OAI21XLTS U247 ( .A0(n59), .A1(n58), .B0(A[2]), .Y(n57) );
  OAI31X1TS U248 ( .A0(n59), .A1(A[2]), .A2(n58), .B0(n57), .Y(n201) );
  INVX2TS U249 ( .A(\mult_x_1/n783 ), .Y(n198) );
  INVX2TS U250 ( .A(B[9]), .Y(n877) );
  INVX2TS U251 ( .A(n323), .Y(n878) );
  OAI22X1TS U252 ( .A0(n152), .A1(n877), .B0(n151), .B1(n878), .Y(n63) );
  OAI22X1TS U253 ( .A0(n153), .A1(n895), .B0(n154), .B1(n893), .Y(n62) );
  OAI21XLTS U254 ( .A0(n63), .A1(n62), .B0(A[2]), .Y(n61) );
  OAI31X1TS U255 ( .A0(n63), .A1(A[2]), .A2(n62), .B0(n61), .Y(n197) );
  INVX2TS U256 ( .A(\mult_x_1/n788 ), .Y(n194) );
  INVX2TS U257 ( .A(B[8]), .Y(n864) );
  INVX2TS U258 ( .A(n326), .Y(n865) );
  OAI22X1TS U259 ( .A0(n152), .A1(n864), .B0(n151), .B1(n865), .Y(n67) );
  OAI22X1TS U260 ( .A0(n153), .A1(n893), .B0(n154), .B1(n877), .Y(n66) );
  OAI21XLTS U261 ( .A0(n67), .A1(n66), .B0(A[2]), .Y(n65) );
  OAI31X1TS U262 ( .A0(n67), .A1(A[2]), .A2(n66), .B0(n65), .Y(n193) );
  INVX2TS U263 ( .A(\mult_x_1/n793 ), .Y(n190) );
  INVX2TS U264 ( .A(B[7]), .Y(n852) );
  INVX2TS U265 ( .A(n329), .Y(n843) );
  OAI22X1TS U266 ( .A0(n152), .A1(n852), .B0(n151), .B1(n843), .Y(n71) );
  OAI22X1TS U267 ( .A0(n153), .A1(n877), .B0(n154), .B1(n864), .Y(n70) );
  OAI21XLTS U268 ( .A0(n71), .A1(n70), .B0(A[2]), .Y(n69) );
  OAI31X1TS U269 ( .A0(n71), .A1(A[2]), .A2(n70), .B0(n69), .Y(n189) );
  INVX2TS U270 ( .A(B[6]), .Y(n885) );
  INVX2TS U271 ( .A(n332), .Y(n847) );
  OAI22X1TS U272 ( .A0(n152), .A1(n885), .B0(n151), .B1(n847), .Y(n75) );
  OAI22X1TS U273 ( .A0(n153), .A1(n864), .B0(n154), .B1(n852), .Y(n74) );
  OAI21XLTS U274 ( .A0(n75), .A1(n74), .B0(A[2]), .Y(n73) );
  OAI31X1TS U275 ( .A0(n75), .A1(A[2]), .A2(n74), .B0(n73), .Y(n186) );
  INVX2TS U276 ( .A(A[6]), .Y(n78) );
  INVX2TS U277 ( .A(A[7]), .Y(n77) );
  OAI22X1TS U278 ( .A0(n78), .A1(A[7]), .B0(n77), .B1(A[6]), .Y(n83) );
  INVX2TS U279 ( .A(A[8]), .Y(n76) );
  AOI22X1TS U280 ( .A0(A[8]), .A1(A[7]), .B0(n77), .B1(n76), .Y(n81) );
  CLKBUFX2TS U281 ( .A(A[5]), .Y(n1036) );
  INVX2TS U282 ( .A(n1036), .Y(n1028) );
  AOI22X1TS U283 ( .A0(n1036), .A1(A[6]), .B0(n78), .B1(n1028), .Y(n87) );
  INVX2TS U284 ( .A(n87), .Y(n82) );
  NAND3BXLTS U285 ( .AN(n83), .B(n81), .C(n82), .Y(n656) );
  OAI21XLTS U286 ( .A0(B[0]), .A1(n817), .B0(n819), .Y(n79) );
  OAI31X1TS U287 ( .A0(B[0]), .A1(n819), .A2(n817), .B0(n79), .Y(n667) );
  OAI22X1TS U288 ( .A0(n928), .A1(n656), .B0(n667), .B1(n80), .Y(n86) );
  NOR2XLTS U289 ( .A(n82), .B(n81), .Y(n964) );
  INVX2TS U290 ( .A(n964), .Y(n820) );
  NAND2X1TS U291 ( .A(n83), .B(n82), .Y(n808) );
  INVX2TS U292 ( .A(n808), .Y(n965) );
  INVX2TS U293 ( .A(n965), .Y(n818) );
  OAI22X1TS U294 ( .A0(n819), .A1(n820), .B0(n817), .B1(n818), .Y(n85) );
  OAI21XLTS U295 ( .A0(n86), .A1(n85), .B0(A[8]), .Y(n84) );
  OAI31X1TS U296 ( .A0(n86), .A1(A[8]), .A2(n85), .B0(n84), .Y(n90) );
  NAND2X1TS U297 ( .A(B[0]), .B(n87), .Y(n122) );
  AOI22X1TS U298 ( .A0(B[1]), .A1(B[0]), .B0(n928), .B1(n817), .Y(n625) );
  INVX2TS U299 ( .A(n625), .Y(n665) );
  OAI222X1TS U300 ( .A0(n80), .A1(n665), .B0(n820), .B1(n817), .C0(n928), .C1(
        n818), .Y(n109) );
  NOR2XLTS U301 ( .A(n76), .B(n109), .Y(n88) );
  NAND2X1TS U302 ( .A(n122), .B(n88), .Y(n89) );
  NOR2XLTS U303 ( .A(n90), .B(n89), .Y(\mult_x_1/n798 ) );
  AO21XLTS U304 ( .A0(n90), .A1(n89), .B0(\mult_x_1/n798 ), .Y(n912) );
  INVX2TS U305 ( .A(A[4]), .Y(n91) );
  OAI22X1TS U306 ( .A0(n1028), .A1(n91), .B0(A[4]), .B1(n1036), .Y(n96) );
  INVX2TS U307 ( .A(A[3]), .Y(n92) );
  AOI22X1TS U308 ( .A0(A[2]), .A1(n92), .B0(A[3]), .B1(n1027), .Y(n150) );
  INVX2TS U309 ( .A(n150), .Y(n135) );
  OAI22X1TS U310 ( .A0(n92), .A1(A[4]), .B0(n91), .B1(A[3]), .Y(n95) );
  NOR2XLTS U311 ( .A(n150), .B(n96), .Y(n100) );
  INVX2TS U312 ( .A(n100), .Y(n1023) );
  INVX2TS U313 ( .A(n350), .Y(n812) );
  OAI22X1TS U314 ( .A0(n819), .A1(n93), .B0(n1023), .B1(n812), .Y(n99) );
  INVX2TS U315 ( .A(B[3]), .Y(n821) );
  NAND2X2TS U316 ( .A(n95), .B(n150), .Y(n904) );
  NAND2X2TS U317 ( .A(n135), .B(n96), .Y(n906) );
  INVX2TS U318 ( .A(B[4]), .Y(n882) );
  OAI22X1TS U319 ( .A0(n821), .A1(n904), .B0(n906), .B1(n882), .Y(n98) );
  OAI21XLTS U320 ( .A0(n99), .A1(n98), .B0(n1036), .Y(n97) );
  OAI31X1TS U321 ( .A0(n99), .A1(n1036), .A2(n98), .B0(n97), .Y(n117) );
  INVX2TS U322 ( .A(n906), .Y(n969) );
  INVX2TS U323 ( .A(n904), .Y(n970) );
  AOI222XLTS U324 ( .A0(B[1]), .A1(n969), .B0(B[0]), .B1(n970), .C0(n625), 
        .C1(n100), .Y(n138) );
  OAI31X1TS U325 ( .A0(n928), .A1(n150), .A2(n1028), .B0(n138), .Y(n136) );
  INVX2TS U326 ( .A(n136), .Y(n104) );
  OAI22X1TS U327 ( .A0(n928), .A1(n93), .B0(n667), .B1(n1023), .Y(n101) );
  AOI21X1TS U328 ( .A0(B[2]), .A1(n969), .B0(n101), .Y(n102) );
  OAI21XLTS U329 ( .A0(n817), .A1(n904), .B0(n102), .Y(n131) );
  NOR2XLTS U330 ( .A(n1028), .B(n131), .Y(n103) );
  NAND2X1TS U331 ( .A(n104), .B(n103), .Y(n130) );
  INVX2TS U332 ( .A(n349), .Y(n816) );
  OAI22X1TS U333 ( .A0(n817), .A1(n93), .B0(n816), .B1(n1023), .Y(n108) );
  OAI22X1TS U334 ( .A0(n821), .A1(n906), .B0(n819), .B1(n904), .Y(n107) );
  OAI21XLTS U335 ( .A0(n108), .A1(n107), .B0(n1036), .Y(n106) );
  OAI31X1TS U336 ( .A0(n108), .A1(n1036), .A2(n107), .B0(n106), .Y(n123) );
  AO21XLTS U337 ( .A0(n122), .A1(n130), .B0(n123), .Y(n116) );
  NOR2XLTS U338 ( .A(n122), .B(n76), .Y(n110) );
  XNOR2X1TS U339 ( .A(n110), .B(n109), .Y(n115) );
  INVX2TS U340 ( .A(n341), .Y(n807) );
  OAI22X1TS U341 ( .A0(n821), .A1(n93), .B0(n1023), .B1(n807), .Y(n114) );
  INVX2TS U342 ( .A(B[5]), .Y(n884) );
  OAI22X1TS U343 ( .A0(n906), .A1(n884), .B0(n904), .B1(n882), .Y(n113) );
  OAI21XLTS U344 ( .A0(n114), .A1(n113), .B0(n1036), .Y(n112) );
  OAI31X1TS U345 ( .A0(n114), .A1(n1036), .A2(n113), .B0(n112), .Y(n910) );
  INVX2TS U346 ( .A(n335), .Y(n851) );
  OAI22X1TS U347 ( .A0(n152), .A1(n884), .B0(n151), .B1(n851), .Y(n121) );
  OAI22X1TS U348 ( .A0(n153), .A1(n852), .B0(n154), .B1(n885), .Y(n120) );
  OAI21XLTS U349 ( .A0(n121), .A1(n120), .B0(A[2]), .Y(n119) );
  OAI31X1TS U350 ( .A0(n121), .A1(A[2]), .A2(n120), .B0(n119), .Y(n181) );
  XOR2XLTS U351 ( .A(n123), .B(n122), .Y(n124) );
  XOR2XLTS U352 ( .A(n130), .B(n124), .Y(n178) );
  INVX2TS U353 ( .A(n338), .Y(n883) );
  OAI22X1TS U354 ( .A0(n152), .A1(n882), .B0(n151), .B1(n883), .Y(n128) );
  OAI22X1TS U355 ( .A0(n153), .A1(n885), .B0(n154), .B1(n884), .Y(n127) );
  OAI21XLTS U356 ( .A0(n128), .A1(n127), .B0(A[2]), .Y(n126) );
  OAI31X1TS U357 ( .A0(n128), .A1(A[2]), .A2(n127), .B0(n126), .Y(n177) );
  NAND3XLTS U358 ( .A(n1036), .B(n136), .C(n131), .Y(n129) );
  OAI211XLTS U359 ( .A0(n1036), .A1(n131), .B0(n130), .C0(n129), .Y(n174) );
  OAI22X1TS U360 ( .A0(n821), .A1(n152), .B0(n151), .B1(n807), .Y(n134) );
  OAI22X1TS U361 ( .A0(n153), .A1(n884), .B0(n154), .B1(n882), .Y(n133) );
  OAI21XLTS U362 ( .A0(n134), .A1(n133), .B0(A[2]), .Y(n132) );
  OAI31X1TS U363 ( .A0(n134), .A1(A[2]), .A2(n133), .B0(n132), .Y(n173) );
  NAND3XLTS U364 ( .A(B[0]), .B(n135), .C(n1036), .Y(n137) );
  OAI21XLTS U365 ( .A0(n138), .A1(n137), .B0(n136), .Y(n170) );
  OAI22X1TS U366 ( .A0(n817), .A1(n152), .B0(n816), .B1(n151), .Y(n141) );
  OAI22X1TS U367 ( .A0(n821), .A1(n153), .B0(n819), .B1(n154), .Y(n140) );
  OAI21XLTS U368 ( .A0(n141), .A1(n140), .B0(n1027), .Y(n139) );
  OAI31X1TS U369 ( .A0(n141), .A1(n1027), .A2(n140), .B0(n139), .Y(n923) );
  NOR2XLTS U370 ( .A(n142), .B(n928), .Y(Product[0]) );
  AOI222XLTS U371 ( .A0(n144), .A1(B[1]), .B0(n143), .B1(B[0]), .C0(n5), .C1(
        n625), .Y(n927) );
  OAI2BB1X1TS U372 ( .A0N(A[2]), .A1N(Product[0]), .B0(n927), .Y(n925) );
  NOR2XLTS U373 ( .A(n1027), .B(n925), .Y(n149) );
  OAI22X1TS U374 ( .A0(n154), .A1(n817), .B0(n151), .B1(n667), .Y(n145) );
  AOI21X1TS U375 ( .A0(n146), .A1(B[0]), .B0(n145), .Y(n147) );
  OAI21XLTS U376 ( .A0(n153), .A1(n819), .B0(n147), .Y(n168) );
  INVX2TS U377 ( .A(n168), .Y(n148) );
  NAND2X1TS U378 ( .A(n149), .B(n148), .Y(n166) );
  OAI21XLTS U379 ( .A0(n928), .A1(n150), .B0(n166), .Y(n924) );
  NAND2X1TS U380 ( .A(n923), .B(n924), .Y(n922) );
  OAI22X1TS U381 ( .A0(n819), .A1(n152), .B0(n151), .B1(n812), .Y(n157) );
  OAI22X1TS U382 ( .A0(n821), .A1(n154), .B0(n153), .B1(n882), .Y(n156) );
  OAI21XLTS U383 ( .A0(n157), .A1(n156), .B0(A[2]), .Y(n155) );
  OAI31X1TS U384 ( .A0(n157), .A1(A[2]), .A2(n156), .B0(n155), .Y(n169) );
  INVX2TS U385 ( .A(n158), .Y(n919) );
  INVX2TS U386 ( .A(n914), .Y(Product[53]) );
  INVX2TS U387 ( .A(n914), .Y(Product[52]) );
  INVX2TS U388 ( .A(n914), .Y(Product[51]) );
  INVX2TS U389 ( .A(A[18]), .Y(n160) );
  INVX2TS U390 ( .A(A[17]), .Y(n1016) );
  AOI22X1TS U391 ( .A0(A[17]), .A1(A[18]), .B0(n160), .B1(n1016), .Y(n465) );
  INVX2TS U392 ( .A(A[19]), .Y(n161) );
  AOI22X1TS U393 ( .A0(A[18]), .A1(n161), .B0(A[19]), .B1(n160), .Y(n163) );
  NOR2XLTS U394 ( .A(n465), .B(n163), .Y(n946) );
  INVX2TS U395 ( .A(n465), .Y(n354) );
  AOI22X1TS U396 ( .A0(A[20]), .A1(A[19]), .B0(n161), .B1(n917), .Y(n355) );
  INVX2TS U397 ( .A(n355), .Y(n162) );
  NOR2XLTS U398 ( .A(n354), .B(n162), .Y(n466) );
  INVX2TS U399 ( .A(n466), .Y(n1012) );
  OAI22X1TS U400 ( .A0(n1012), .A1(n1009), .B0(n1011), .B1(n1001), .Y(n165) );
  OAI21XLTS U401 ( .A0(n946), .A1(n165), .B0(n917), .Y(n164) );
  OAI31X1TS U402 ( .A0(n946), .A1(n917), .A2(n165), .B0(n164), .Y(
        \mult_x_1/n1057 ) );
  INVX2TS U403 ( .A(A[14]), .Y(n1035) );
  INVX2TS U404 ( .A(\mult_x_1/n363 ), .Y(\mult_x_1/n373 ) );
  INVX2TS U405 ( .A(A[21]), .Y(n284) );
  AOI22X1TS U406 ( .A0(A[20]), .A1(n284), .B0(A[21]), .B1(n917), .Y(n286) );
  NOR2XLTS U407 ( .A(n286), .B(n928), .Y(\mult_x_1/n705 ) );
  OAI21XLTS U408 ( .A0(n168), .A1(A[2]), .B0(n166), .Y(n167) );
  AOI31XLTS U409 ( .A0(n168), .A1(A[2]), .A2(n925), .B0(n167), .Y(Product[2])
         );
  INVX2TS U410 ( .A(n171), .Y(Product[4]) );
  INVX2TS U411 ( .A(n175), .Y(Product[5]) );
  INVX2TS U412 ( .A(n179), .Y(Product[6]) );
  INVX2TS U413 ( .A(n183), .Y(Product[7]) );
  INVX2TS U414 ( .A(n187), .Y(Product[8]) );
  INVX2TS U415 ( .A(n191), .Y(Product[9]) );
  INVX2TS U416 ( .A(n195), .Y(Product[10]) );
  INVX2TS U417 ( .A(n199), .Y(Product[11]) );
  INVX2TS U418 ( .A(n203), .Y(Product[12]) );
  INVX2TS U419 ( .A(n207), .Y(Product[13]) );
  INVX2TS U420 ( .A(n211), .Y(Product[14]) );
  NOR2XLTS U421 ( .A(A[2]), .B(n1036), .Y(n242) );
  INVX2TS U422 ( .A(n242), .Y(n1026) );
  NOR2XLTS U423 ( .A(n1026), .B(A[8]), .Y(n1025) );
  NOR2XLTS U424 ( .A(\mult_x_1/n448 ), .B(n1025), .Y(n283) );
  INVX2TS U425 ( .A(n212), .Y(\mult_x_1/n413 ) );
  INVX2TS U426 ( .A(n216), .Y(Product[15]) );
  INVX2TS U427 ( .A(n220), .Y(Product[16]) );
  INVX2TS U428 ( .A(n221), .Y(\mult_x_1/n414 ) );
  INVX2TS U429 ( .A(n225), .Y(Product[17]) );
  INVX2TS U430 ( .A(n229), .Y(Product[18]) );
  INVX2TS U431 ( .A(n233), .Y(Product[19]) );
  INVX2TS U432 ( .A(n237), .Y(Product[20]) );
  INVX2TS U433 ( .A(n241), .Y(Product[21]) );
  AOI211XLTS U434 ( .A0(n1036), .A1(A[2]), .B0(n242), .C0(n1030), .Y(
        \mult_x_1/n463 ) );
  NOR2XLTS U435 ( .A(n242), .B(\mult_x_1/n463 ), .Y(\mult_x_1/n464 ) );
  INVX2TS U436 ( .A(n246), .Y(Product[22]) );
  INVX2TS U437 ( .A(n250), .Y(Product[23]) );
  INVX2TS U438 ( .A(n254), .Y(Product[24]) );
  INVX2TS U439 ( .A(n258), .Y(Product[25]) );
  INVX2TS U440 ( .A(n261), .Y(Product[26]) );
  INVX2TS U441 ( .A(n264), .Y(Product[27]) );
  INVX2TS U442 ( .A(n267), .Y(Product[28]) );
  INVX2TS U443 ( .A(n270), .Y(Product[29]) );
  INVX2TS U444 ( .A(n273), .Y(Product[30]) );
  INVX2TS U445 ( .A(n276), .Y(Product[31]) );
  INVX2TS U446 ( .A(n279), .Y(Product[32]) );
  INVX2TS U447 ( .A(n282), .Y(Product[33]) );
  INVX2TS U448 ( .A(n283), .Y(n301) );
  AOI21X1TS U449 ( .A0(\mult_x_1/n448 ), .A1(n1025), .B0(n283), .Y(n298) );
  NOR3XLTS U450 ( .A(A[20]), .B(A[21]), .C(A[22]), .Y(n346) );
  CLKBUFX2TS U451 ( .A(n346), .Y(n1008) );
  INVX2TS U452 ( .A(A[22]), .Y(n285) );
  OAI33XLTS U453 ( .A0(A[20]), .A1(A[21]), .A2(n285), .B0(n917), .B1(n284), 
        .B2(A[22]), .Y(n295) );
  CLKBUFX2TS U454 ( .A(n295), .Y(n999) );
  AOI22X1TS U455 ( .A0(n1008), .A1(B[18]), .B0(n999), .B1(B[19]), .Y(n289) );
  NOR2X2TS U456 ( .A(n286), .B(A[22]), .Y(n1010) );
  NOR2X2TS U457 ( .A(n286), .B(n285), .Y(n983) );
  AOI22X1TS U458 ( .A0(n1010), .A1(n287), .B0(n983), .B1(B[20]), .Y(n288) );
  NAND2X1TS U459 ( .A(n289), .B(n288), .Y(n297) );
  INVX2TS U460 ( .A(n290), .Y(\mult_x_1/n424 ) );
  INVX2TS U461 ( .A(n294), .Y(Product[34]) );
  INVX2TS U462 ( .A(n1010), .Y(n1006) );
  INVX2TS U463 ( .A(n295), .Y(n1005) );
  OAI22X1TS U464 ( .A0(n967), .A1(n1006), .B0(n1005), .B1(n1001), .Y(n296) );
  AOI211XLTS U465 ( .A0(n1008), .A1(B[21]), .B0(n983), .C0(n296), .Y(
        \mult_x_1/n1023 ) );
  INVX2TS U466 ( .A(n299), .Y(\mult_x_1/n438 ) );
  INVX2TS U467 ( .A(n302), .Y(\mult_x_1/n425 ) );
  INVX2TS U468 ( .A(n306), .Y(Product[35]) );
  INVX2TS U469 ( .A(n310), .Y(Product[36]) );
  INVX2TS U470 ( .A(n983), .Y(n1002) );
  AOI22X1TS U471 ( .A0(n1008), .A1(B[11]), .B0(n999), .B1(B[12]), .Y(n311) );
  OAI21XLTS U472 ( .A0(n1002), .A1(n1030), .B0(n311), .Y(n312) );
  AOI21X1TS U473 ( .A0(n1010), .A1(n313), .B0(n312), .Y(n921) );
  INVX2TS U474 ( .A(n318), .Y(Product[37]) );
  AOI22X1TS U475 ( .A0(n1008), .A1(B[10]), .B0(n999), .B1(B[11]), .Y(n322) );
  AOI22X1TS U476 ( .A0(n1010), .A1(n320), .B0(n983), .B1(B[12]), .Y(n321) );
  NAND2X1TS U477 ( .A(n322), .B(n321), .Y(n370) );
  AOI22X1TS U478 ( .A0(n1008), .A1(B[9]), .B0(n999), .B1(B[10]), .Y(n325) );
  AOI22X1TS U479 ( .A0(n1010), .A1(n323), .B0(n983), .B1(B[11]), .Y(n324) );
  NAND2X1TS U480 ( .A(n325), .B(n324), .Y(n391) );
  AOI22X1TS U481 ( .A0(n1008), .A1(B[8]), .B0(n999), .B1(B[9]), .Y(n328) );
  AOI22X1TS U482 ( .A0(n1010), .A1(n326), .B0(n983), .B1(B[10]), .Y(n327) );
  NAND2X1TS U483 ( .A(n328), .B(n327), .Y(n388) );
  AOI22X1TS U484 ( .A0(n1008), .A1(B[7]), .B0(n999), .B1(B[8]), .Y(n331) );
  AOI22X1TS U485 ( .A0(n1010), .A1(n329), .B0(n983), .B1(B[9]), .Y(n330) );
  NAND2X1TS U486 ( .A(n331), .B(n330), .Y(n385) );
  AOI22X1TS U487 ( .A0(n1008), .A1(B[6]), .B0(n999), .B1(B[7]), .Y(n334) );
  AOI22X1TS U488 ( .A0(n1010), .A1(n332), .B0(n983), .B1(B[8]), .Y(n333) );
  NAND2X1TS U489 ( .A(n334), .B(n333), .Y(n382) );
  AOI22X1TS U490 ( .A0(n1008), .A1(B[5]), .B0(n999), .B1(B[6]), .Y(n337) );
  AOI22X1TS U491 ( .A0(n1010), .A1(n335), .B0(n983), .B1(B[7]), .Y(n336) );
  NAND2X1TS U492 ( .A(n337), .B(n336), .Y(n379) );
  AOI22X1TS U493 ( .A0(n1008), .A1(B[4]), .B0(n999), .B1(B[5]), .Y(n340) );
  AOI22X1TS U494 ( .A0(n1010), .A1(n338), .B0(n983), .B1(B[6]), .Y(n339) );
  NAND2X1TS U495 ( .A(n340), .B(n339), .Y(n373) );
  AOI22X1TS U496 ( .A0(B[3]), .A1(n1008), .B0(n999), .B1(B[4]), .Y(n343) );
  AOI22X1TS U497 ( .A0(n1010), .A1(n341), .B0(n983), .B1(B[5]), .Y(n342) );
  NAND2X1TS U498 ( .A(n343), .B(n342), .Y(n376) );
  INVX2TS U499 ( .A(\mult_x_1/n705 ), .Y(n934) );
  AOI222XLTS U500 ( .A0(B[1]), .A1(n983), .B0(B[0]), .B1(n999), .C0(n625), 
        .C1(n1010), .Y(n935) );
  NAND2X1TS U501 ( .A(n934), .B(n935), .Y(n933) );
  AOI22X1TS U502 ( .A0(B[1]), .A1(n999), .B0(B[0]), .B1(n346), .Y(n345) );
  NAND2X1TS U503 ( .A(B[2]), .B(n983), .Y(n344) );
  OAI211XLTS U504 ( .A0(n1006), .A1(n667), .B0(n345), .C0(n344), .Y(n932) );
  NOR2XLTS U505 ( .A(n933), .B(n932), .Y(n931) );
  AOI22X1TS U506 ( .A0(B[2]), .A1(n999), .B0(B[1]), .B1(n346), .Y(n347) );
  OAI21XLTS U507 ( .A0(n821), .A1(n1002), .B0(n347), .Y(n348) );
  AOI21X1TS U508 ( .A0(n349), .A1(n1010), .B0(n348), .Y(n929) );
  OAI21XLTS U509 ( .A0(B[0]), .A1(n931), .B0(n929), .Y(n394) );
  AOI22X1TS U510 ( .A0(B[3]), .A1(n999), .B0(B[2]), .B1(n1008), .Y(n352) );
  AOI22X1TS U511 ( .A0(n1010), .A1(n350), .B0(n983), .B1(B[4]), .Y(n351) );
  NAND2X1TS U512 ( .A(n352), .B(n351), .Y(n393) );
  INVX2TS U513 ( .A(n353), .Y(\mult_x_1/n546 ) );
  OAI22X1TS U514 ( .A0(n1012), .A1(n835), .B0(n1011), .B1(\mult_x_1/n404 ), 
        .Y(n358) );
  NOR2XLTS U515 ( .A(n355), .B(n354), .Y(n945) );
  INVX2TS U516 ( .A(n945), .Y(n475) );
  INVX2TS U517 ( .A(n946), .Y(n474) );
  OAI22X1TS U518 ( .A0(n475), .A1(n1001), .B0(n474), .B1(n996), .Y(n357) );
  OAI21XLTS U519 ( .A0(n358), .A1(n357), .B0(n917), .Y(n356) );
  OAI31X1TS U520 ( .A0(n358), .A1(n917), .A2(n357), .B0(n356), .Y(
        \mult_x_1/n1059 ) );
  OAI22X1TS U521 ( .A0(n1012), .A1(n831), .B0(n1011), .B1(n992), .Y(n361) );
  OAI22X1TS U522 ( .A0(n475), .A1(n996), .B0(n474), .B1(\mult_x_1/n404 ), .Y(
        n360) );
  OAI21XLTS U523 ( .A0(n361), .A1(n360), .B0(n917), .Y(n359) );
  OAI31X1TS U524 ( .A0(n361), .A1(n917), .A2(n360), .B0(n359), .Y(
        \mult_x_1/n1060 ) );
  INVX2TS U525 ( .A(n365), .Y(Product[38]) );
  OAI22X1TS U526 ( .A0(n1012), .A1(n889), .B0(n1011), .B1(n988), .Y(n368) );
  OAI22X1TS U527 ( .A0(n475), .A1(\mult_x_1/n404 ), .B0(n474), .B1(n992), .Y(
        n367) );
  OAI21XLTS U528 ( .A0(n368), .A1(n367), .B0(n917), .Y(n366) );
  OAI31X1TS U529 ( .A0(n368), .A1(n917), .A2(n367), .B0(n366), .Y(
        \mult_x_1/n1061 ) );
  INVX2TS U530 ( .A(n371), .Y(\mult_x_1/n547 ) );
  INVX2TS U531 ( .A(n374), .Y(\mult_x_1/n631 ) );
  INVX2TS U532 ( .A(n377), .Y(\mult_x_1/n644 ) );
  INVX2TS U533 ( .A(n380), .Y(\mult_x_1/n617 ) );
  INVX2TS U534 ( .A(n383), .Y(\mult_x_1/n603 ) );
  INVX2TS U535 ( .A(n386), .Y(\mult_x_1/n589 ) );
  INVX2TS U536 ( .A(n389), .Y(\mult_x_1/n575 ) );
  INVX2TS U537 ( .A(n392), .Y(\mult_x_1/n561 ) );
  INVX2TS U538 ( .A(n395), .Y(\mult_x_1/n657 ) );
  OAI22X1TS U539 ( .A0(n1012), .A1(n856), .B0(n1011), .B1(n905), .Y(n398) );
  OAI22X1TS U540 ( .A0(n475), .A1(n992), .B0(n474), .B1(n988), .Y(n397) );
  OAI21XLTS U541 ( .A0(n398), .A1(n397), .B0(n917), .Y(n396) );
  OAI31X1TS U542 ( .A0(n398), .A1(n917), .A2(n397), .B0(n396), .Y(
        \mult_x_1/n1062 ) );
  INVX2TS U543 ( .A(n402), .Y(Product[39]) );
  XNOR2X1TS U544 ( .A(A[15]), .B(A[16]), .Y(n405) );
  AOI2BB2XLTS U545 ( .B0(A[15]), .B1(n1035), .A0N(n1035), .A1N(A[15]), .Y(n495) );
  INVX2TS U546 ( .A(n495), .Y(n403) );
  NOR2XLTS U547 ( .A(n405), .B(n403), .Y(n950) );
  AOI2BB2XLTS U548 ( .B0(A[17]), .B1(A[16]), .A0N(A[16]), .A1N(A[17]), .Y(n451) );
  NAND3XLTS U549 ( .A(n451), .B(n495), .C(n405), .Y(n1014) );
  OAI22X1TS U550 ( .A0(n404), .A1(n1009), .B0(n1014), .B1(n1001), .Y(n407) );
  OAI21XLTS U551 ( .A0(n950), .A1(n407), .B0(n1016), .Y(n406) );
  OAI31X1TS U552 ( .A0(n950), .A1(n1016), .A2(n407), .B0(n406), .Y(
        \mult_x_1/n1092 ) );
  OAI22X1TS U553 ( .A0(n1012), .A1(n869), .B0(n1011), .B1(n903), .Y(n410) );
  OAI22X1TS U554 ( .A0(n475), .A1(n988), .B0(n474), .B1(n905), .Y(n409) );
  OAI21XLTS U555 ( .A0(n410), .A1(n409), .B0(n917), .Y(n408) );
  OAI31X1TS U556 ( .A0(n410), .A1(n917), .A2(n409), .B0(n408), .Y(
        \mult_x_1/n1063 ) );
  OAI22X1TS U557 ( .A0(n1012), .A1(n985), .B0(n1011), .B1(n977), .Y(n413) );
  OAI22X1TS U558 ( .A0(n475), .A1(n905), .B0(n474), .B1(n903), .Y(n412) );
  OAI21XLTS U559 ( .A0(n413), .A1(n412), .B0(n917), .Y(n411) );
  OAI31X1TS U560 ( .A0(n413), .A1(n917), .A2(n412), .B0(n411), .Y(
        \mult_x_1/n1064 ) );
  OAI22X1TS U561 ( .A0(n1012), .A1(n981), .B0(n1011), .B1(n973), .Y(n416) );
  OAI22X1TS U562 ( .A0(n475), .A1(n903), .B0(n474), .B1(n977), .Y(n415) );
  OAI21XLTS U563 ( .A0(n416), .A1(n415), .B0(n917), .Y(n414) );
  OAI31X1TS U564 ( .A0(n416), .A1(n917), .A2(n415), .B0(n414), .Y(
        \mult_x_1/n1065 ) );
  INVX2TS U565 ( .A(n420), .Y(Product[40]) );
  OAI22X1TS U566 ( .A0(n1012), .A1(n860), .B0(n1011), .B1(n1030), .Y(n423) );
  OAI22X1TS U567 ( .A0(n475), .A1(n977), .B0(n474), .B1(n973), .Y(n422) );
  OAI21XLTS U568 ( .A0(n423), .A1(n422), .B0(n917), .Y(n421) );
  OAI31X1TS U569 ( .A0(n423), .A1(n917), .A2(n422), .B0(n421), .Y(
        \mult_x_1/n1066 ) );
  OAI22X1TS U570 ( .A0(n1012), .A1(n847), .B0(n1011), .B1(n885), .Y(n426) );
  OAI22X1TS U571 ( .A0(n475), .A1(n864), .B0(n474), .B1(n852), .Y(n425) );
  OAI21XLTS U572 ( .A0(n426), .A1(n425), .B0(n917), .Y(n424) );
  OAI31X1TS U573 ( .A0(n426), .A1(n917), .A2(n425), .B0(n424), .Y(
        \mult_x_1/n1073 ) );
  OAI22X1TS U574 ( .A0(n1012), .A1(n851), .B0(n1011), .B1(n884), .Y(n429) );
  OAI22X1TS U575 ( .A0(n475), .A1(n852), .B0(n474), .B1(n885), .Y(n428) );
  OAI21XLTS U576 ( .A0(n429), .A1(n428), .B0(n917), .Y(n427) );
  OAI31X1TS U577 ( .A0(n429), .A1(n917), .A2(n428), .B0(n427), .Y(
        \mult_x_1/n1074 ) );
  OAI22X1TS U578 ( .A0(n1012), .A1(n865), .B0(n1011), .B1(n864), .Y(n432) );
  OAI22X1TS U579 ( .A0(n475), .A1(n893), .B0(n474), .B1(n877), .Y(n431) );
  OAI21XLTS U580 ( .A0(n432), .A1(n431), .B0(n917), .Y(n430) );
  OAI31X1TS U581 ( .A0(n432), .A1(n917), .A2(n431), .B0(n430), .Y(
        \mult_x_1/n1071 ) );
  OAI22X1TS U582 ( .A0(n1012), .A1(n843), .B0(n1011), .B1(n852), .Y(n435) );
  OAI22X1TS U583 ( .A0(n475), .A1(n877), .B0(n474), .B1(n864), .Y(n434) );
  OAI21XLTS U584 ( .A0(n435), .A1(n434), .B0(n917), .Y(n433) );
  OAI31X1TS U585 ( .A0(n435), .A1(n917), .A2(n434), .B0(n433), .Y(
        \mult_x_1/n1072 ) );
  OAI22X1TS U586 ( .A0(n1012), .A1(n883), .B0(n1011), .B1(n882), .Y(n438) );
  OAI22X1TS U587 ( .A0(n475), .A1(n885), .B0(n474), .B1(n884), .Y(n437) );
  OAI21XLTS U588 ( .A0(n438), .A1(n437), .B0(n917), .Y(n436) );
  OAI31X1TS U589 ( .A0(n438), .A1(n917), .A2(n437), .B0(n436), .Y(
        \mult_x_1/n1075 ) );
  OAI22X1TS U590 ( .A0(n1012), .A1(n894), .B0(n1011), .B1(n893), .Y(n441) );
  OAI22X1TS U591 ( .A0(n475), .A1(n896), .B0(n474), .B1(n895), .Y(n440) );
  OAI21XLTS U592 ( .A0(n441), .A1(n440), .B0(n917), .Y(n439) );
  OAI31X1TS U593 ( .A0(n441), .A1(n917), .A2(n440), .B0(n439), .Y(
        \mult_x_1/n1069 ) );
  OAI22X1TS U594 ( .A0(n1012), .A1(n878), .B0(n1011), .B1(n877), .Y(n444) );
  OAI22X1TS U595 ( .A0(n475), .A1(n895), .B0(n474), .B1(n893), .Y(n443) );
  OAI21XLTS U596 ( .A0(n444), .A1(n443), .B0(n917), .Y(n442) );
  OAI31X1TS U597 ( .A0(n444), .A1(n917), .A2(n443), .B0(n442), .Y(
        \mult_x_1/n1070 ) );
  OAI22X1TS U598 ( .A0(n1012), .A1(n839), .B0(n1011), .B1(n895), .Y(n447) );
  OAI22X1TS U599 ( .A0(n475), .A1(n1030), .B0(n474), .B1(n896), .Y(n446) );
  OAI21XLTS U600 ( .A0(n447), .A1(n446), .B0(n917), .Y(n445) );
  OAI31X1TS U601 ( .A0(n447), .A1(n917), .A2(n446), .B0(n445), .Y(
        \mult_x_1/n1068 ) );
  OAI22X1TS U602 ( .A0(n1012), .A1(n873), .B0(n1011), .B1(n896), .Y(n450) );
  OAI22X1TS U603 ( .A0(n475), .A1(n973), .B0(n474), .B1(n1030), .Y(n449) );
  OAI21XLTS U604 ( .A0(n450), .A1(n449), .B0(n917), .Y(n448) );
  OAI31X1TS U605 ( .A0(n450), .A1(n917), .A2(n449), .B0(n448), .Y(
        \mult_x_1/n1067 ) );
  CLKBUFX2TS U606 ( .A(n1014), .Y(n568) );
  OAI22X1TS U607 ( .A0(n404), .A1(n835), .B0(n568), .B1(\mult_x_1/n404 ), .Y(
        n454) );
  NOR2XLTS U608 ( .A(n495), .B(n451), .Y(n949) );
  INVX2TS U609 ( .A(n949), .Y(n570) );
  INVX2TS U610 ( .A(n950), .Y(n569) );
  OAI22X1TS U611 ( .A0(n570), .A1(n1001), .B0(n569), .B1(n996), .Y(n453) );
  OAI21XLTS U612 ( .A0(n454), .A1(n453), .B0(n1016), .Y(n452) );
  OAI31X1TS U613 ( .A0(n454), .A1(n1016), .A2(n453), .B0(n452), .Y(
        \mult_x_1/n1094 ) );
  OAI22X1TS U614 ( .A0(n821), .A1(n1011), .B0(n1012), .B1(n807), .Y(n457) );
  OAI22X1TS U615 ( .A0(n475), .A1(n884), .B0(n474), .B1(n882), .Y(n456) );
  OAI21XLTS U616 ( .A0(n457), .A1(n456), .B0(n917), .Y(n455) );
  OAI31X1TS U617 ( .A0(n457), .A1(n917), .A2(n456), .B0(n455), .Y(
        \mult_x_1/n1076 ) );
  OAI22X1TS U618 ( .A0(n819), .A1(n1011), .B0(n1012), .B1(n812), .Y(n460) );
  OAI22X1TS U619 ( .A0(n821), .A1(n474), .B0(n475), .B1(n882), .Y(n459) );
  OAI21XLTS U620 ( .A0(n460), .A1(n459), .B0(n917), .Y(n458) );
  OAI31X1TS U621 ( .A0(n460), .A1(n917), .A2(n459), .B0(n458), .Y(
        \mult_x_1/n1077 ) );
  INVX2TS U622 ( .A(n464), .Y(Product[41]) );
  NAND2X1TS U623 ( .A(B[0]), .B(n465), .Y(n514) );
  AOI222XLTS U624 ( .A0(B[1]), .A1(n945), .B0(B[0]), .B1(n946), .C0(n625), 
        .C1(n466), .Y(n515) );
  OAI21XLTS U625 ( .A0(n514), .A1(n917), .B0(n515), .Y(n513) );
  INVX2TS U626 ( .A(n513), .Y(n557) );
  NAND2X1TS U627 ( .A(A[20]), .B(n557), .Y(n470) );
  AOI2BB2XLTS U628 ( .B0(B[2]), .B1(n945), .A0N(n928), .A1N(n1011), .Y(n467)
         );
  OAI21XLTS U629 ( .A0(n667), .A1(n1012), .B0(n467), .Y(n468) );
  AOI21X1TS U630 ( .A0(B[1]), .A1(n946), .B0(n468), .Y(n556) );
  INVX2TS U631 ( .A(n556), .Y(n469) );
  NOR2XLTS U632 ( .A(n470), .B(n469), .Y(\mult_x_1/n714 ) );
  OAI22X1TS U633 ( .A0(n404), .A1(n831), .B0(n568), .B1(n992), .Y(n473) );
  OAI22X1TS U634 ( .A0(n570), .A1(n996), .B0(n569), .B1(\mult_x_1/n404 ), .Y(
        n472) );
  OAI21XLTS U635 ( .A0(n473), .A1(n472), .B0(n1016), .Y(n471) );
  OAI31X1TS U636 ( .A0(n473), .A1(n1016), .A2(n472), .B0(n471), .Y(
        \mult_x_1/n1095 ) );
  OAI22X1TS U637 ( .A0(n817), .A1(n1011), .B0(n816), .B1(n1012), .Y(n478) );
  OAI22X1TS U638 ( .A0(n821), .A1(n475), .B0(n819), .B1(n474), .Y(n477) );
  OAI21XLTS U639 ( .A0(n478), .A1(n477), .B0(n917), .Y(n476) );
  OAI31X1TS U640 ( .A0(n478), .A1(n917), .A2(n477), .B0(n476), .Y(
        \mult_x_1/n1078 ) );
  OAI22X1TS U641 ( .A0(n404), .A1(n889), .B0(n568), .B1(n988), .Y(n481) );
  OAI22X1TS U642 ( .A0(n570), .A1(\mult_x_1/n404 ), .B0(n569), .B1(n992), .Y(
        n480) );
  OAI21XLTS U643 ( .A0(n481), .A1(n480), .B0(n1016), .Y(n479) );
  OAI31X1TS U644 ( .A0(n481), .A1(n1016), .A2(n480), .B0(n479), .Y(
        \mult_x_1/n1096 ) );
  OAI22X1TS U645 ( .A0(n404), .A1(n856), .B0(n568), .B1(n905), .Y(n484) );
  OAI22X1TS U646 ( .A0(n570), .A1(n992), .B0(n569), .B1(n988), .Y(n483) );
  OAI21XLTS U647 ( .A0(n484), .A1(n483), .B0(n1016), .Y(n482) );
  OAI31X1TS U648 ( .A0(n484), .A1(n1016), .A2(n483), .B0(n482), .Y(
        \mult_x_1/n1097 ) );
  INVX2TS U649 ( .A(n488), .Y(Product[42]) );
  INVX2TS U650 ( .A(A[12]), .Y(n489) );
  INVX2TS U651 ( .A(A[11]), .Y(n957) );
  AOI22X1TS U652 ( .A0(A[11]), .A1(A[12]), .B0(n489), .B1(n957), .Y(n623) );
  INVX2TS U653 ( .A(A[13]), .Y(n490) );
  AOI22X1TS U654 ( .A0(A[12]), .A1(n490), .B0(A[13]), .B1(n489), .Y(n492) );
  NOR2XLTS U655 ( .A(n623), .B(n492), .Y(n954) );
  INVX2TS U656 ( .A(n623), .Y(n523) );
  AOI22X1TS U657 ( .A0(A[14]), .A1(A[13]), .B0(n490), .B1(n1035), .Y(n524) );
  INVX2TS U658 ( .A(n524), .Y(n491) );
  NOR2XLTS U659 ( .A(n523), .B(n491), .Y(n624) );
  INVX2TS U660 ( .A(n624), .Y(n1018) );
  OAI22X1TS U661 ( .A0(n1018), .A1(n1009), .B0(n1017), .B1(n1001), .Y(n494) );
  OAI21XLTS U662 ( .A0(n954), .A1(n494), .B0(n1035), .Y(n493) );
  OAI31X1TS U663 ( .A0(n954), .A1(n1035), .A2(n494), .B0(n493), .Y(
        \mult_x_1/n1127 ) );
  NOR2XLTS U664 ( .A(n928), .B(n495), .Y(\mult_x_1/n759 ) );
  OAI222X1TS U665 ( .A0(n404), .A1(n665), .B0(n570), .B1(n817), .C0(n569), 
        .C1(n928), .Y(n496) );
  AOI21X1TS U666 ( .A0(A[17]), .A1(\mult_x_1/n759 ), .B0(n496), .Y(n937) );
  AOI31XLTS U667 ( .A0(A[17]), .A1(\mult_x_1/n759 ), .A2(n496), .B0(n937), .Y(
        \mult_x_1/n751 ) );
  NAND2X1TS U668 ( .A(A[17]), .B(n937), .Y(n500) );
  OAI22X1TS U669 ( .A0(n928), .A1(n1014), .B0(n667), .B1(n404), .Y(n498) );
  OAI22X1TS U670 ( .A0(n819), .A1(n570), .B0(n817), .B1(n569), .Y(n497) );
  NOR2XLTS U671 ( .A(n498), .B(n497), .Y(n939) );
  INVX2TS U672 ( .A(n939), .Y(n499) );
  OR2X1TS U673 ( .A(n500), .B(n499), .Y(n936) );
  OAI22X1TS U674 ( .A0(n817), .A1(n568), .B0(n816), .B1(n404), .Y(n503) );
  OAI22X1TS U675 ( .A0(n821), .A1(n570), .B0(n819), .B1(n569), .Y(n502) );
  OAI21XLTS U676 ( .A0(n503), .A1(n502), .B0(A[17]), .Y(n501) );
  OAI31X1TS U677 ( .A0(n503), .A1(A[17]), .A2(n502), .B0(n501), .Y(n512) );
  XNOR2X1TS U678 ( .A(n936), .B(n512), .Y(n504) );
  XOR2XLTS U679 ( .A(n514), .B(n504), .Y(\mult_x_1/n733 ) );
  INVX2TS U680 ( .A(n508), .Y(Product[43]) );
  OAI22X1TS U681 ( .A0(n819), .A1(n568), .B0(n404), .B1(n812), .Y(n511) );
  OAI22X1TS U682 ( .A0(n821), .A1(n569), .B0(n570), .B1(n882), .Y(n510) );
  OAI21XLTS U683 ( .A0(n511), .A1(n510), .B0(A[17]), .Y(n509) );
  OAI31X1TS U684 ( .A0(n511), .A1(A[17]), .A2(n510), .B0(n509), .Y(n560) );
  AO21XLTS U685 ( .A0(n936), .A1(n514), .B0(n512), .Y(n559) );
  OAI31X1TS U686 ( .A0(n515), .A1(n917), .A2(n514), .B0(n513), .Y(n558) );
  INVX2TS U687 ( .A(n516), .Y(\mult_x_1/n723 ) );
  OAI22X1TS U688 ( .A0(n404), .A1(n869), .B0(n568), .B1(n903), .Y(n519) );
  OAI22X1TS U689 ( .A0(n570), .A1(n988), .B0(n569), .B1(n905), .Y(n518) );
  OAI21XLTS U690 ( .A0(n519), .A1(n518), .B0(n1016), .Y(n517) );
  OAI31X1TS U691 ( .A0(n519), .A1(n1016), .A2(n518), .B0(n517), .Y(
        \mult_x_1/n1098 ) );
  OAI22X1TS U692 ( .A0(n404), .A1(n839), .B0(n568), .B1(n895), .Y(n522) );
  OAI22X1TS U693 ( .A0(n570), .A1(n1030), .B0(n569), .B1(n896), .Y(n521) );
  OAI21XLTS U694 ( .A0(n522), .A1(n521), .B0(n1016), .Y(n520) );
  OAI31X1TS U695 ( .A0(n522), .A1(n1016), .A2(n521), .B0(n520), .Y(
        \mult_x_1/n1103 ) );
  OAI22X1TS U696 ( .A0(n1018), .A1(n835), .B0(n1017), .B1(\mult_x_1/n404 ), 
        .Y(n527) );
  NOR2XLTS U697 ( .A(n524), .B(n523), .Y(n953) );
  INVX2TS U698 ( .A(n953), .Y(n643) );
  INVX2TS U699 ( .A(n954), .Y(n642) );
  OAI22X1TS U700 ( .A0(n643), .A1(n1001), .B0(n642), .B1(n996), .Y(n526) );
  OAI21XLTS U701 ( .A0(n527), .A1(n526), .B0(n1035), .Y(n525) );
  OAI31X1TS U702 ( .A0(n527), .A1(n1035), .A2(n526), .B0(n525), .Y(
        \mult_x_1/n1129 ) );
  OAI22X1TS U703 ( .A0(n404), .A1(n847), .B0(n568), .B1(n885), .Y(n530) );
  OAI22X1TS U704 ( .A0(n570), .A1(n864), .B0(n569), .B1(n852), .Y(n529) );
  OAI21XLTS U705 ( .A0(n530), .A1(n529), .B0(n1016), .Y(n528) );
  OAI31X1TS U706 ( .A0(n530), .A1(n1016), .A2(n529), .B0(n528), .Y(
        \mult_x_1/n1108 ) );
  OAI22X1TS U707 ( .A0(n404), .A1(n878), .B0(n568), .B1(n877), .Y(n533) );
  OAI22X1TS U708 ( .A0(n570), .A1(n895), .B0(n569), .B1(n893), .Y(n532) );
  OAI21XLTS U709 ( .A0(n533), .A1(n532), .B0(n1016), .Y(n531) );
  OAI31X1TS U710 ( .A0(n533), .A1(n1016), .A2(n532), .B0(n531), .Y(
        \mult_x_1/n1105 ) );
  OAI22X1TS U711 ( .A0(n404), .A1(n851), .B0(n568), .B1(n884), .Y(n536) );
  OAI22X1TS U712 ( .A0(n570), .A1(n852), .B0(n569), .B1(n885), .Y(n535) );
  OAI21XLTS U713 ( .A0(n536), .A1(n535), .B0(n1016), .Y(n534) );
  OAI31X1TS U714 ( .A0(n536), .A1(n1016), .A2(n535), .B0(n534), .Y(
        \mult_x_1/n1109 ) );
  OAI22X1TS U715 ( .A0(n404), .A1(n843), .B0(n568), .B1(n852), .Y(n539) );
  OAI22X1TS U716 ( .A0(n570), .A1(n877), .B0(n569), .B1(n864), .Y(n538) );
  OAI21XLTS U717 ( .A0(n539), .A1(n538), .B0(n1016), .Y(n537) );
  OAI31X1TS U718 ( .A0(n539), .A1(n1016), .A2(n538), .B0(n537), .Y(
        \mult_x_1/n1107 ) );
  OAI22X1TS U719 ( .A0(n404), .A1(n894), .B0(n568), .B1(n893), .Y(n542) );
  OAI22X1TS U720 ( .A0(n570), .A1(n896), .B0(n569), .B1(n895), .Y(n541) );
  OAI21XLTS U721 ( .A0(n542), .A1(n541), .B0(n1016), .Y(n540) );
  OAI31X1TS U722 ( .A0(n542), .A1(n1016), .A2(n541), .B0(n540), .Y(
        \mult_x_1/n1104 ) );
  OAI22X1TS U723 ( .A0(n404), .A1(n883), .B0(n568), .B1(n882), .Y(n545) );
  OAI22X1TS U724 ( .A0(n570), .A1(n885), .B0(n569), .B1(n884), .Y(n544) );
  OAI21XLTS U725 ( .A0(n545), .A1(n544), .B0(n1016), .Y(n543) );
  OAI31X1TS U726 ( .A0(n545), .A1(n1016), .A2(n544), .B0(n543), .Y(
        \mult_x_1/n1110 ) );
  OAI22X1TS U727 ( .A0(n404), .A1(n865), .B0(n568), .B1(n864), .Y(n548) );
  OAI22X1TS U728 ( .A0(n570), .A1(n893), .B0(n569), .B1(n877), .Y(n547) );
  OAI21XLTS U729 ( .A0(n548), .A1(n547), .B0(n1016), .Y(n546) );
  OAI31X1TS U730 ( .A0(n548), .A1(n1016), .A2(n547), .B0(n546), .Y(
        \mult_x_1/n1106 ) );
  OAI22X1TS U731 ( .A0(n404), .A1(n873), .B0(n568), .B1(n896), .Y(n551) );
  OAI22X1TS U732 ( .A0(n570), .A1(n973), .B0(n569), .B1(n1030), .Y(n550) );
  OAI21XLTS U733 ( .A0(n551), .A1(n550), .B0(n1016), .Y(n549) );
  OAI31X1TS U734 ( .A0(n551), .A1(n1016), .A2(n550), .B0(n549), .Y(
        \mult_x_1/n1102 ) );
  OAI22X1TS U735 ( .A0(n404), .A1(n860), .B0(n568), .B1(n1030), .Y(n554) );
  OAI22X1TS U736 ( .A0(n570), .A1(n977), .B0(n569), .B1(n973), .Y(n553) );
  OAI21XLTS U737 ( .A0(n554), .A1(n553), .B0(n1016), .Y(n552) );
  OAI31X1TS U738 ( .A0(n554), .A1(n1016), .A2(n553), .B0(n552), .Y(
        \mult_x_1/n1101 ) );
  OAI21XLTS U739 ( .A0(n557), .A1(n917), .B0(n556), .Y(n555) );
  OAI31X1TS U740 ( .A0(n557), .A1(n556), .A2(n917), .B0(n555), .Y(n576) );
  OAI22X1TS U741 ( .A0(n821), .A1(n568), .B0(n404), .B1(n807), .Y(n563) );
  OAI22X1TS U742 ( .A0(n570), .A1(n884), .B0(n569), .B1(n882), .Y(n562) );
  OAI21XLTS U743 ( .A0(n563), .A1(n562), .B0(A[17]), .Y(n561) );
  OAI31X1TS U744 ( .A0(n563), .A1(A[17]), .A2(n562), .B0(n561), .Y(n574) );
  INVX2TS U745 ( .A(n564), .Y(\mult_x_1/n712 ) );
  OAI22X1TS U746 ( .A0(n404), .A1(n981), .B0(n568), .B1(n973), .Y(n567) );
  OAI22X1TS U747 ( .A0(n570), .A1(n903), .B0(n569), .B1(n977), .Y(n566) );
  OAI21XLTS U748 ( .A0(n567), .A1(n566), .B0(n1016), .Y(n565) );
  OAI31X1TS U749 ( .A0(n567), .A1(n1016), .A2(n566), .B0(n565), .Y(
        \mult_x_1/n1100 ) );
  OAI22X1TS U750 ( .A0(n404), .A1(n985), .B0(n568), .B1(n977), .Y(n573) );
  OAI22X1TS U751 ( .A0(n570), .A1(n905), .B0(n569), .B1(n903), .Y(n572) );
  OAI21XLTS U752 ( .A0(n573), .A1(n572), .B0(n1016), .Y(n571) );
  OAI31X1TS U753 ( .A0(n573), .A1(n1016), .A2(n572), .B0(n571), .Y(
        \mult_x_1/n1099 ) );
  INVX2TS U754 ( .A(n577), .Y(\mult_x_1/n713 ) );
  OAI22X1TS U755 ( .A0(n1018), .A1(n831), .B0(n1017), .B1(n992), .Y(n580) );
  OAI22X1TS U756 ( .A0(n643), .A1(n996), .B0(n642), .B1(\mult_x_1/n404 ), .Y(
        n579) );
  OAI21XLTS U757 ( .A0(n580), .A1(n579), .B0(n1035), .Y(n578) );
  OAI31X1TS U758 ( .A0(n580), .A1(n1035), .A2(n579), .B0(n578), .Y(
        \mult_x_1/n1130 ) );
  OAI22X1TS U759 ( .A0(n1018), .A1(n860), .B0(n1017), .B1(n1030), .Y(n583) );
  OAI22X1TS U760 ( .A0(n643), .A1(n977), .B0(n642), .B1(n973), .Y(n582) );
  OAI21XLTS U761 ( .A0(n583), .A1(n582), .B0(n1035), .Y(n581) );
  OAI31X1TS U762 ( .A0(n583), .A1(n1035), .A2(n582), .B0(n581), .Y(
        \mult_x_1/n1136 ) );
  OAI22X1TS U763 ( .A0(n1018), .A1(n839), .B0(n1017), .B1(n895), .Y(n586) );
  OAI22X1TS U764 ( .A0(n643), .A1(n1030), .B0(n642), .B1(n896), .Y(n585) );
  OAI21XLTS U765 ( .A0(n586), .A1(n585), .B0(n1035), .Y(n584) );
  OAI31X1TS U766 ( .A0(n586), .A1(n1035), .A2(n585), .B0(n584), .Y(
        \mult_x_1/n1138 ) );
  OAI22X1TS U767 ( .A0(n1018), .A1(n873), .B0(n1017), .B1(n896), .Y(n589) );
  OAI22X1TS U768 ( .A0(n643), .A1(n973), .B0(n642), .B1(n1030), .Y(n588) );
  OAI21XLTS U769 ( .A0(n589), .A1(n588), .B0(n1035), .Y(n587) );
  OAI31X1TS U770 ( .A0(n589), .A1(n1035), .A2(n588), .B0(n587), .Y(
        \mult_x_1/n1137 ) );
  OAI22X1TS U771 ( .A0(n1018), .A1(n843), .B0(n1017), .B1(n852), .Y(n592) );
  OAI22X1TS U772 ( .A0(n643), .A1(n877), .B0(n642), .B1(n864), .Y(n591) );
  OAI21XLTS U773 ( .A0(n592), .A1(n591), .B0(n1035), .Y(n590) );
  OAI31X1TS U774 ( .A0(n592), .A1(n1035), .A2(n591), .B0(n590), .Y(
        \mult_x_1/n1142 ) );
  OAI22X1TS U775 ( .A0(n1018), .A1(n851), .B0(n1017), .B1(n884), .Y(n595) );
  OAI22X1TS U776 ( .A0(n643), .A1(n852), .B0(n642), .B1(n885), .Y(n594) );
  OAI21XLTS U777 ( .A0(n595), .A1(n594), .B0(n1035), .Y(n593) );
  OAI31X1TS U778 ( .A0(n595), .A1(n1035), .A2(n594), .B0(n593), .Y(
        \mult_x_1/n1144 ) );
  OAI22X1TS U779 ( .A0(n1018), .A1(n847), .B0(n1017), .B1(n885), .Y(n598) );
  OAI22X1TS U780 ( .A0(n643), .A1(n864), .B0(n642), .B1(n852), .Y(n597) );
  OAI21XLTS U781 ( .A0(n598), .A1(n597), .B0(n1035), .Y(n596) );
  OAI31X1TS U782 ( .A0(n598), .A1(n1035), .A2(n597), .B0(n596), .Y(
        \mult_x_1/n1143 ) );
  OAI22X1TS U783 ( .A0(n1018), .A1(n865), .B0(n1017), .B1(n864), .Y(n601) );
  OAI22X1TS U784 ( .A0(n643), .A1(n893), .B0(n642), .B1(n877), .Y(n600) );
  OAI21XLTS U785 ( .A0(n601), .A1(n600), .B0(n1035), .Y(n599) );
  OAI31X1TS U786 ( .A0(n601), .A1(n1035), .A2(n600), .B0(n599), .Y(
        \mult_x_1/n1141 ) );
  OAI22X1TS U787 ( .A0(n1018), .A1(n883), .B0(n1017), .B1(n882), .Y(n604) );
  OAI22X1TS U788 ( .A0(n643), .A1(n885), .B0(n642), .B1(n884), .Y(n603) );
  OAI21XLTS U789 ( .A0(n604), .A1(n603), .B0(n1035), .Y(n602) );
  OAI31X1TS U790 ( .A0(n604), .A1(n1035), .A2(n603), .B0(n602), .Y(
        \mult_x_1/n1145 ) );
  OAI22X1TS U791 ( .A0(n1018), .A1(n878), .B0(n1017), .B1(n877), .Y(n607) );
  OAI22X1TS U792 ( .A0(n643), .A1(n895), .B0(n642), .B1(n893), .Y(n606) );
  OAI21XLTS U793 ( .A0(n607), .A1(n606), .B0(n1035), .Y(n605) );
  OAI31X1TS U794 ( .A0(n607), .A1(n1035), .A2(n606), .B0(n605), .Y(
        \mult_x_1/n1140 ) );
  OAI22X1TS U795 ( .A0(n1018), .A1(n894), .B0(n1017), .B1(n893), .Y(n610) );
  OAI22X1TS U796 ( .A0(n643), .A1(n896), .B0(n642), .B1(n895), .Y(n609) );
  OAI21XLTS U797 ( .A0(n610), .A1(n609), .B0(n1035), .Y(n608) );
  OAI31X1TS U798 ( .A0(n610), .A1(n1035), .A2(n609), .B0(n608), .Y(
        \mult_x_1/n1139 ) );
  OAI22X1TS U799 ( .A0(n1018), .A1(n869), .B0(n1017), .B1(n903), .Y(n613) );
  OAI22X1TS U800 ( .A0(n643), .A1(n988), .B0(n642), .B1(n905), .Y(n612) );
  OAI21XLTS U801 ( .A0(n613), .A1(n612), .B0(n1035), .Y(n611) );
  OAI31X1TS U802 ( .A0(n613), .A1(n1035), .A2(n612), .B0(n611), .Y(
        \mult_x_1/n1133 ) );
  OAI22X1TS U803 ( .A0(n1018), .A1(n981), .B0(n1017), .B1(n973), .Y(n616) );
  OAI22X1TS U804 ( .A0(n643), .A1(n903), .B0(n642), .B1(n977), .Y(n615) );
  OAI21XLTS U805 ( .A0(n616), .A1(n615), .B0(n1035), .Y(n614) );
  OAI31X1TS U806 ( .A0(n616), .A1(n1035), .A2(n615), .B0(n614), .Y(
        \mult_x_1/n1135 ) );
  OAI22X1TS U807 ( .A0(n1018), .A1(n985), .B0(n1017), .B1(n977), .Y(n619) );
  OAI22X1TS U808 ( .A0(n643), .A1(n905), .B0(n642), .B1(n903), .Y(n618) );
  OAI21XLTS U809 ( .A0(n619), .A1(n618), .B0(n1035), .Y(n617) );
  OAI31X1TS U810 ( .A0(n619), .A1(n1035), .A2(n618), .B0(n617), .Y(
        \mult_x_1/n1134 ) );
  OAI22X1TS U811 ( .A0(n1018), .A1(n856), .B0(n1017), .B1(n905), .Y(n622) );
  OAI22X1TS U812 ( .A0(n643), .A1(n992), .B0(n642), .B1(n988), .Y(n621) );
  OAI21XLTS U813 ( .A0(n622), .A1(n621), .B0(n1035), .Y(n620) );
  OAI31X1TS U814 ( .A0(n622), .A1(n1035), .A2(n621), .B0(n620), .Y(
        \mult_x_1/n1132 ) );
  NAND2X1TS U815 ( .A(B[0]), .B(n623), .Y(n680) );
  AOI222XLTS U816 ( .A0(B[1]), .A1(n953), .B0(B[0]), .B1(n954), .C0(n625), 
        .C1(n624), .Y(n681) );
  OAI21XLTS U817 ( .A0(n1035), .A1(n680), .B0(n681), .Y(n683) );
  AOI2BB2XLTS U818 ( .B0(B[2]), .B1(n953), .A0N(n928), .A1N(n1017), .Y(n626)
         );
  OAI21XLTS U819 ( .A0(n667), .A1(n1018), .B0(n626), .Y(n627) );
  AOI21X1TS U820 ( .A0(B[1]), .A1(n954), .B0(n627), .Y(n685) );
  NAND2X1TS U821 ( .A(A[14]), .B(n685), .Y(n628) );
  NOR2XLTS U822 ( .A(n683), .B(n628), .Y(\mult_x_1/n765 ) );
  OAI22X1TS U823 ( .A0(n1018), .A1(n889), .B0(n1017), .B1(n988), .Y(n631) );
  OAI22X1TS U824 ( .A0(n643), .A1(\mult_x_1/n404 ), .B0(n642), .B1(n992), .Y(
        n630) );
  OAI21XLTS U825 ( .A0(n631), .A1(n630), .B0(n1035), .Y(n629) );
  OAI31X1TS U826 ( .A0(n631), .A1(n1035), .A2(n630), .B0(n629), .Y(
        \mult_x_1/n1131 ) );
  INVX2TS U827 ( .A(n635), .Y(Product[44]) );
  OAI22X1TS U828 ( .A0(n821), .A1(n1017), .B0(n1018), .B1(n807), .Y(n638) );
  OAI22X1TS U829 ( .A0(n643), .A1(n884), .B0(n642), .B1(n882), .Y(n637) );
  OAI21XLTS U830 ( .A0(n638), .A1(n637), .B0(n1035), .Y(n636) );
  OAI31X1TS U831 ( .A0(n638), .A1(n1035), .A2(n637), .B0(n636), .Y(
        \mult_x_1/n1146 ) );
  OAI22X1TS U832 ( .A0(n819), .A1(n1017), .B0(n1018), .B1(n812), .Y(n641) );
  OAI22X1TS U833 ( .A0(n821), .A1(n642), .B0(n643), .B1(n882), .Y(n640) );
  OAI21XLTS U834 ( .A0(n641), .A1(n640), .B0(n1035), .Y(n639) );
  OAI31X1TS U835 ( .A0(n641), .A1(n1035), .A2(n640), .B0(n639), .Y(
        \mult_x_1/n1147 ) );
  OAI22X1TS U836 ( .A0(n817), .A1(n1017), .B0(n816), .B1(n1018), .Y(n646) );
  OAI22X1TS U837 ( .A0(n821), .A1(n643), .B0(n819), .B1(n642), .Y(n645) );
  OAI21XLTS U838 ( .A0(n646), .A1(n645), .B0(n1035), .Y(n644) );
  OAI31X1TS U839 ( .A0(n646), .A1(n1035), .A2(n645), .B0(n644), .Y(
        \mult_x_1/n1148 ) );
  INVX2TS U840 ( .A(n650), .Y(Product[45]) );
  XNOR2X1TS U841 ( .A(A[10]), .B(A[9]), .Y(n653) );
  AOI2BB2XLTS U842 ( .B0(A[9]), .B1(n76), .A0N(n76), .A1N(A[9]), .Y(n664) );
  INVX2TS U843 ( .A(n664), .Y(n651) );
  NOR2XLTS U844 ( .A(n653), .B(n651), .Y(n961) );
  AOI2BB2XLTS U845 ( .B0(A[11]), .B1(A[10]), .A0N(A[10]), .A1N(A[11]), .Y(n663) );
  NAND3XLTS U846 ( .A(n663), .B(n664), .C(n653), .Y(n958) );
  OAI22X1TS U847 ( .A0(n652), .A1(n1009), .B0(n958), .B1(n1001), .Y(n655) );
  OAI21XLTS U848 ( .A0(n961), .A1(n655), .B0(n957), .Y(n654) );
  OAI31X1TS U849 ( .A0(n961), .A1(n957), .A2(n655), .B0(n654), .Y(
        \mult_x_1/n1162 ) );
  CLKBUFX2TS U850 ( .A(n656), .Y(n1020) );
  OAI22X1TS U851 ( .A0(n80), .A1(n1009), .B0(n1020), .B1(n1001), .Y(n658) );
  OAI21XLTS U852 ( .A0(n965), .A1(n658), .B0(n76), .Y(n657) );
  OAI31X1TS U853 ( .A0(n965), .A1(n76), .A2(n658), .B0(n657), .Y(
        \mult_x_1/n1197 ) );
  INVX2TS U854 ( .A(n662), .Y(Product[46]) );
  NOR2XLTS U855 ( .A(n928), .B(n664), .Y(\mult_x_1/n795 ) );
  NOR2XLTS U856 ( .A(n664), .B(n663), .Y(n960) );
  INVX2TS U857 ( .A(n960), .Y(n742) );
  INVX2TS U858 ( .A(n961), .Y(n744) );
  OAI222X1TS U859 ( .A0(n652), .A1(n665), .B0(n742), .B1(n817), .C0(n744), 
        .C1(n928), .Y(n666) );
  AOI21X1TS U860 ( .A0(A[11]), .A1(\mult_x_1/n795 ), .B0(n666), .Y(n941) );
  AOI31XLTS U861 ( .A0(A[11]), .A1(\mult_x_1/n795 ), .A2(n666), .B0(n941), .Y(
        \mult_x_1/n790 ) );
  NAND2X1TS U862 ( .A(A[11]), .B(n941), .Y(n671) );
  OAI22X1TS U863 ( .A0(n819), .A1(n742), .B0(n667), .B1(n652), .Y(n669) );
  OAI22X1TS U864 ( .A0(n817), .A1(n744), .B0(n928), .B1(n958), .Y(n668) );
  NOR2XLTS U865 ( .A(n669), .B(n668), .Y(n943) );
  INVX2TS U866 ( .A(n943), .Y(n670) );
  OR2X1TS U867 ( .A(n671), .B(n670), .Y(n940) );
  OAI22X1TS U868 ( .A0(n821), .A1(n742), .B0(n816), .B1(n652), .Y(n674) );
  CLKBUFX2TS U869 ( .A(n958), .Y(n743) );
  OAI22X1TS U870 ( .A0(n819), .A1(n744), .B0(n817), .B1(n743), .Y(n673) );
  OAI21XLTS U871 ( .A0(n674), .A1(n673), .B0(A[11]), .Y(n672) );
  OAI31X1TS U872 ( .A0(n674), .A1(A[11]), .A2(n673), .B0(n672), .Y(n679) );
  XNOR2X1TS U873 ( .A(n940), .B(n679), .Y(n675) );
  XOR2XLTS U874 ( .A(n680), .B(n675), .Y(\mult_x_1/n778 ) );
  OAI22X1TS U875 ( .A0(n742), .A1(n882), .B0(n652), .B1(n812), .Y(n678) );
  OAI22X1TS U876 ( .A0(n821), .A1(n744), .B0(n819), .B1(n743), .Y(n677) );
  OAI21XLTS U877 ( .A0(n678), .A1(n677), .B0(A[11]), .Y(n676) );
  OAI31X1TS U878 ( .A0(n678), .A1(A[11]), .A2(n677), .B0(n676), .Y(n689) );
  AO21XLTS U879 ( .A0(n940), .A1(n680), .B0(n679), .Y(n688) );
  OAI31X1TS U880 ( .A0(n681), .A1(n680), .A2(n1035), .B0(n683), .Y(n687) );
  INVX2TS U881 ( .A(n682), .Y(\mult_x_1/n771 ) );
  INVX2TS U882 ( .A(n683), .Y(n686) );
  OAI21XLTS U883 ( .A0(n686), .A1(n1035), .B0(n685), .Y(n684) );
  OAI31X1TS U884 ( .A0(n686), .A1(n685), .A2(n1035), .B0(n684), .Y(n750) );
  OAI22X1TS U885 ( .A0(n742), .A1(n884), .B0(n652), .B1(n807), .Y(n692) );
  OAI22X1TS U886 ( .A0(n821), .A1(n743), .B0(n744), .B1(n882), .Y(n691) );
  OAI21XLTS U887 ( .A0(n692), .A1(n691), .B0(A[11]), .Y(n690) );
  OAI31X1TS U888 ( .A0(n692), .A1(A[11]), .A2(n691), .B0(n690), .Y(n748) );
  INVX2TS U889 ( .A(n693), .Y(\mult_x_1/n763 ) );
  OAI22X1TS U890 ( .A0(n742), .A1(n992), .B0(n652), .B1(n856), .Y(n696) );
  OAI22X1TS U891 ( .A0(n744), .A1(n988), .B0(n743), .B1(n905), .Y(n695) );
  OAI21XLTS U892 ( .A0(n696), .A1(n695), .B0(n957), .Y(n694) );
  OAI31X1TS U893 ( .A0(n696), .A1(n957), .A2(n695), .B0(n694), .Y(
        \mult_x_1/n1167 ) );
  OAI22X1TS U894 ( .A0(n742), .A1(n852), .B0(n652), .B1(n851), .Y(n699) );
  OAI22X1TS U895 ( .A0(n744), .A1(n885), .B0(n743), .B1(n884), .Y(n698) );
  OAI21XLTS U896 ( .A0(n699), .A1(n698), .B0(n957), .Y(n697) );
  OAI31X1TS U897 ( .A0(n699), .A1(n957), .A2(n698), .B0(n697), .Y(
        \mult_x_1/n1179 ) );
  OAI22X1TS U898 ( .A0(n742), .A1(n1030), .B0(n652), .B1(n839), .Y(n702) );
  OAI22X1TS U899 ( .A0(n744), .A1(n896), .B0(n743), .B1(n895), .Y(n701) );
  OAI21XLTS U900 ( .A0(n702), .A1(n701), .B0(n957), .Y(n700) );
  OAI31X1TS U901 ( .A0(n702), .A1(n957), .A2(n701), .B0(n700), .Y(
        \mult_x_1/n1173 ) );
  OAI22X1TS U902 ( .A0(n742), .A1(n973), .B0(n652), .B1(n873), .Y(n705) );
  OAI22X1TS U903 ( .A0(n744), .A1(n1030), .B0(n743), .B1(n896), .Y(n704) );
  OAI21XLTS U904 ( .A0(n705), .A1(n704), .B0(n957), .Y(n703) );
  OAI31X1TS U905 ( .A0(n705), .A1(n957), .A2(n704), .B0(n703), .Y(
        \mult_x_1/n1172 ) );
  OAI22X1TS U906 ( .A0(n742), .A1(n977), .B0(n652), .B1(n860), .Y(n708) );
  OAI22X1TS U907 ( .A0(n744), .A1(n973), .B0(n743), .B1(n1030), .Y(n707) );
  OAI21XLTS U908 ( .A0(n708), .A1(n707), .B0(n957), .Y(n706) );
  OAI31X1TS U909 ( .A0(n708), .A1(n957), .A2(n707), .B0(n706), .Y(
        \mult_x_1/n1171 ) );
  OAI22X1TS U910 ( .A0(n742), .A1(n895), .B0(n652), .B1(n878), .Y(n711) );
  OAI22X1TS U911 ( .A0(n744), .A1(n893), .B0(n743), .B1(n877), .Y(n710) );
  OAI21XLTS U912 ( .A0(n711), .A1(n710), .B0(n957), .Y(n709) );
  OAI31X1TS U913 ( .A0(n711), .A1(n957), .A2(n710), .B0(n709), .Y(
        \mult_x_1/n1175 ) );
  OAI22X1TS U914 ( .A0(n742), .A1(n864), .B0(n652), .B1(n847), .Y(n714) );
  OAI22X1TS U915 ( .A0(n744), .A1(n852), .B0(n743), .B1(n885), .Y(n713) );
  OAI21XLTS U916 ( .A0(n714), .A1(n713), .B0(n957), .Y(n712) );
  OAI31X1TS U917 ( .A0(n714), .A1(n957), .A2(n713), .B0(n712), .Y(
        \mult_x_1/n1178 ) );
  OAI22X1TS U918 ( .A0(n742), .A1(n896), .B0(n652), .B1(n894), .Y(n717) );
  OAI22X1TS U919 ( .A0(n744), .A1(n895), .B0(n743), .B1(n893), .Y(n716) );
  OAI21XLTS U920 ( .A0(n717), .A1(n716), .B0(n957), .Y(n715) );
  OAI31X1TS U921 ( .A0(n717), .A1(n957), .A2(n716), .B0(n715), .Y(
        \mult_x_1/n1174 ) );
  OAI22X1TS U922 ( .A0(n742), .A1(n885), .B0(n652), .B1(n883), .Y(n720) );
  OAI22X1TS U923 ( .A0(n744), .A1(n884), .B0(n743), .B1(n882), .Y(n719) );
  OAI21XLTS U924 ( .A0(n720), .A1(n719), .B0(n957), .Y(n718) );
  OAI31X1TS U925 ( .A0(n720), .A1(n957), .A2(n719), .B0(n718), .Y(
        \mult_x_1/n1180 ) );
  OAI22X1TS U926 ( .A0(n742), .A1(n988), .B0(n652), .B1(n869), .Y(n723) );
  OAI22X1TS U927 ( .A0(n744), .A1(n905), .B0(n743), .B1(n903), .Y(n722) );
  OAI21XLTS U928 ( .A0(n723), .A1(n722), .B0(n957), .Y(n721) );
  OAI31X1TS U929 ( .A0(n723), .A1(n957), .A2(n722), .B0(n721), .Y(
        \mult_x_1/n1168 ) );
  OAI22X1TS U930 ( .A0(n742), .A1(n1001), .B0(n652), .B1(n835), .Y(n726) );
  OAI22X1TS U931 ( .A0(n744), .A1(n996), .B0(n958), .B1(\mult_x_1/n404 ), .Y(
        n725) );
  OAI21XLTS U932 ( .A0(n726), .A1(n725), .B0(n957), .Y(n724) );
  OAI31X1TS U933 ( .A0(n726), .A1(n957), .A2(n725), .B0(n724), .Y(
        \mult_x_1/n1164 ) );
  OAI22X1TS U934 ( .A0(n742), .A1(n996), .B0(n652), .B1(n831), .Y(n729) );
  OAI22X1TS U935 ( .A0(n744), .A1(\mult_x_1/n404 ), .B0(n958), .B1(n992), .Y(
        n728) );
  OAI21XLTS U936 ( .A0(n729), .A1(n728), .B0(n957), .Y(n727) );
  OAI31X1TS U937 ( .A0(n729), .A1(n957), .A2(n728), .B0(n727), .Y(
        \mult_x_1/n1165 ) );
  OAI22X1TS U938 ( .A0(n742), .A1(n893), .B0(n652), .B1(n865), .Y(n732) );
  OAI22X1TS U939 ( .A0(n744), .A1(n877), .B0(n743), .B1(n864), .Y(n731) );
  OAI21XLTS U940 ( .A0(n732), .A1(n731), .B0(n957), .Y(n730) );
  OAI31X1TS U941 ( .A0(n732), .A1(n957), .A2(n731), .B0(n730), .Y(
        \mult_x_1/n1176 ) );
  OAI22X1TS U942 ( .A0(n742), .A1(n877), .B0(n652), .B1(n843), .Y(n735) );
  OAI22X1TS U943 ( .A0(n744), .A1(n864), .B0(n743), .B1(n852), .Y(n734) );
  OAI21XLTS U944 ( .A0(n735), .A1(n734), .B0(n957), .Y(n733) );
  OAI31X1TS U945 ( .A0(n735), .A1(n957), .A2(n734), .B0(n733), .Y(
        \mult_x_1/n1177 ) );
  OAI22X1TS U946 ( .A0(n742), .A1(\mult_x_1/n404 ), .B0(n652), .B1(n889), .Y(
        n738) );
  OAI22X1TS U947 ( .A0(n744), .A1(n992), .B0(n743), .B1(n988), .Y(n737) );
  OAI21XLTS U948 ( .A0(n738), .A1(n737), .B0(n957), .Y(n736) );
  OAI31X1TS U949 ( .A0(n738), .A1(n957), .A2(n737), .B0(n736), .Y(
        \mult_x_1/n1166 ) );
  OAI22X1TS U950 ( .A0(n742), .A1(n905), .B0(n652), .B1(n985), .Y(n741) );
  OAI22X1TS U951 ( .A0(n744), .A1(n903), .B0(n743), .B1(n977), .Y(n740) );
  OAI21XLTS U952 ( .A0(n741), .A1(n740), .B0(n957), .Y(n739) );
  OAI31X1TS U953 ( .A0(n741), .A1(n957), .A2(n740), .B0(n739), .Y(
        \mult_x_1/n1169 ) );
  OAI22X1TS U954 ( .A0(n742), .A1(n903), .B0(n652), .B1(n981), .Y(n747) );
  OAI22X1TS U955 ( .A0(n744), .A1(n977), .B0(n743), .B1(n973), .Y(n746) );
  OAI21XLTS U956 ( .A0(n747), .A1(n746), .B0(n957), .Y(n745) );
  OAI31X1TS U957 ( .A0(n747), .A1(n957), .A2(n746), .B0(n745), .Y(
        \mult_x_1/n1170 ) );
  INVX2TS U958 ( .A(n751), .Y(\mult_x_1/n764 ) );
  OAI22X1TS U959 ( .A0(n80), .A1(n839), .B0(n1020), .B1(n895), .Y(n754) );
  OAI22X1TS U960 ( .A0(n808), .A1(n896), .B0(n820), .B1(n1030), .Y(n753) );
  OAI21XLTS U961 ( .A0(n754), .A1(n753), .B0(n76), .Y(n752) );
  OAI31X1TS U962 ( .A0(n754), .A1(n76), .A2(n753), .B0(n752), .Y(
        \mult_x_1/n1208 ) );
  OAI22X1TS U963 ( .A0(n80), .A1(n860), .B0(n1020), .B1(n1030), .Y(n757) );
  OAI22X1TS U964 ( .A0(n808), .A1(n973), .B0(n820), .B1(n977), .Y(n756) );
  OAI21XLTS U965 ( .A0(n757), .A1(n756), .B0(n76), .Y(n755) );
  OAI31X1TS U966 ( .A0(n757), .A1(n76), .A2(n756), .B0(n755), .Y(
        \mult_x_1/n1206 ) );
  OAI22X1TS U967 ( .A0(n80), .A1(n873), .B0(n1020), .B1(n896), .Y(n760) );
  OAI22X1TS U968 ( .A0(n818), .A1(n1030), .B0(n820), .B1(n973), .Y(n759) );
  OAI21XLTS U969 ( .A0(n760), .A1(n759), .B0(n76), .Y(n758) );
  OAI31X1TS U970 ( .A0(n760), .A1(n76), .A2(n759), .B0(n758), .Y(
        \mult_x_1/n1207 ) );
  OAI22X1TS U971 ( .A0(n80), .A1(n856), .B0(n1020), .B1(n905), .Y(n763) );
  OAI22X1TS U972 ( .A0(n818), .A1(n988), .B0(n820), .B1(n992), .Y(n762) );
  OAI21XLTS U973 ( .A0(n763), .A1(n762), .B0(n76), .Y(n761) );
  OAI31X1TS U974 ( .A0(n763), .A1(n76), .A2(n762), .B0(n761), .Y(
        \mult_x_1/n1202 ) );
  OAI22X1TS U975 ( .A0(n80), .A1(n869), .B0(n1020), .B1(n903), .Y(n766) );
  OAI22X1TS U976 ( .A0(n808), .A1(n905), .B0(n820), .B1(n988), .Y(n765) );
  OAI21XLTS U977 ( .A0(n766), .A1(n765), .B0(n76), .Y(n764) );
  OAI31X1TS U978 ( .A0(n766), .A1(n76), .A2(n765), .B0(n764), .Y(
        \mult_x_1/n1203 ) );
  OAI22X1TS U979 ( .A0(n80), .A1(n831), .B0(n1020), .B1(n992), .Y(n769) );
  OAI22X1TS U980 ( .A0(n808), .A1(\mult_x_1/n404 ), .B0(n820), .B1(n996), .Y(
        n768) );
  OAI21XLTS U981 ( .A0(n769), .A1(n768), .B0(n76), .Y(n767) );
  OAI31X1TS U982 ( .A0(n769), .A1(n76), .A2(n768), .B0(n767), .Y(
        \mult_x_1/n1200 ) );
  OAI22X1TS U983 ( .A0(n80), .A1(n894), .B0(n1020), .B1(n893), .Y(n772) );
  OAI22X1TS U984 ( .A0(n808), .A1(n895), .B0(n820), .B1(n896), .Y(n771) );
  OAI21XLTS U985 ( .A0(n772), .A1(n771), .B0(n76), .Y(n770) );
  OAI31X1TS U986 ( .A0(n772), .A1(n76), .A2(n771), .B0(n770), .Y(
        \mult_x_1/n1209 ) );
  OAI22X1TS U987 ( .A0(n80), .A1(n865), .B0(n1020), .B1(n864), .Y(n775) );
  OAI22X1TS U988 ( .A0(n808), .A1(n877), .B0(n820), .B1(n893), .Y(n774) );
  OAI21XLTS U989 ( .A0(n775), .A1(n774), .B0(n76), .Y(n773) );
  OAI31X1TS U990 ( .A0(n775), .A1(n76), .A2(n774), .B0(n773), .Y(
        \mult_x_1/n1211 ) );
  OAI22X1TS U991 ( .A0(n80), .A1(n835), .B0(n1020), .B1(\mult_x_1/n404 ), .Y(
        n778) );
  OAI22X1TS U992 ( .A0(n818), .A1(n996), .B0(n820), .B1(n1001), .Y(n777) );
  OAI21XLTS U993 ( .A0(n778), .A1(n777), .B0(n76), .Y(n776) );
  OAI31X1TS U994 ( .A0(n778), .A1(n76), .A2(n777), .B0(n776), .Y(
        \mult_x_1/n1199 ) );
  OAI22X1TS U995 ( .A0(n80), .A1(n878), .B0(n1020), .B1(n877), .Y(n781) );
  OAI22X1TS U996 ( .A0(n808), .A1(n893), .B0(n820), .B1(n895), .Y(n780) );
  OAI21XLTS U997 ( .A0(n781), .A1(n780), .B0(n76), .Y(n779) );
  OAI31X1TS U998 ( .A0(n781), .A1(n76), .A2(n780), .B0(n779), .Y(
        \mult_x_1/n1210 ) );
  OAI22X1TS U999 ( .A0(n80), .A1(n843), .B0(n1020), .B1(n852), .Y(n784) );
  OAI22X1TS U1000 ( .A0(n818), .A1(n864), .B0(n820), .B1(n877), .Y(n783) );
  OAI21XLTS U1001 ( .A0(n784), .A1(n783), .B0(n76), .Y(n782) );
  OAI31X1TS U1002 ( .A0(n784), .A1(n76), .A2(n783), .B0(n782), .Y(
        \mult_x_1/n1212 ) );
  OAI22X1TS U1003 ( .A0(n80), .A1(n847), .B0(n1020), .B1(n885), .Y(n787) );
  OAI22X1TS U1004 ( .A0(n808), .A1(n852), .B0(n820), .B1(n864), .Y(n786) );
  OAI21XLTS U1005 ( .A0(n787), .A1(n786), .B0(n76), .Y(n785) );
  OAI31X1TS U1006 ( .A0(n787), .A1(n76), .A2(n786), .B0(n785), .Y(
        \mult_x_1/n1213 ) );
  OAI22X1TS U1007 ( .A0(n80), .A1(n851), .B0(n1020), .B1(n884), .Y(n790) );
  OAI22X1TS U1008 ( .A0(n808), .A1(n885), .B0(n820), .B1(n852), .Y(n789) );
  OAI21XLTS U1009 ( .A0(n790), .A1(n789), .B0(n76), .Y(n788) );
  OAI31X1TS U1010 ( .A0(n790), .A1(n76), .A2(n789), .B0(n788), .Y(
        \mult_x_1/n1214 ) );
  OAI22X1TS U1011 ( .A0(n80), .A1(n889), .B0(n1020), .B1(n988), .Y(n793) );
  OAI22X1TS U1012 ( .A0(n808), .A1(n992), .B0(n820), .B1(\mult_x_1/n404 ), .Y(
        n792) );
  OAI21XLTS U1013 ( .A0(n793), .A1(n792), .B0(n76), .Y(n791) );
  OAI31X1TS U1014 ( .A0(n793), .A1(n76), .A2(n792), .B0(n791), .Y(
        \mult_x_1/n1201 ) );
  OAI22X1TS U1015 ( .A0(n80), .A1(n883), .B0(n1020), .B1(n882), .Y(n796) );
  OAI22X1TS U1016 ( .A0(n808), .A1(n884), .B0(n820), .B1(n885), .Y(n795) );
  OAI21XLTS U1017 ( .A0(n796), .A1(n795), .B0(n76), .Y(n794) );
  OAI31X1TS U1018 ( .A0(n796), .A1(n76), .A2(n795), .B0(n794), .Y(
        \mult_x_1/n1215 ) );
  OAI22X1TS U1019 ( .A0(n80), .A1(n981), .B0(n1020), .B1(n973), .Y(n799) );
  OAI22X1TS U1020 ( .A0(n818), .A1(n977), .B0(n820), .B1(n903), .Y(n798) );
  OAI21XLTS U1021 ( .A0(n799), .A1(n798), .B0(n76), .Y(n797) );
  OAI31X1TS U1022 ( .A0(n799), .A1(n76), .A2(n798), .B0(n797), .Y(
        \mult_x_1/n1205 ) );
  OAI22X1TS U1023 ( .A0(n80), .A1(n985), .B0(n1020), .B1(n977), .Y(n802) );
  OAI22X1TS U1024 ( .A0(n818), .A1(n903), .B0(n820), .B1(n905), .Y(n801) );
  OAI21XLTS U1025 ( .A0(n802), .A1(n801), .B0(n76), .Y(n800) );
  OAI31X1TS U1026 ( .A0(n802), .A1(n76), .A2(n801), .B0(n800), .Y(
        \mult_x_1/n1204 ) );
  INVX2TS U1027 ( .A(n806), .Y(Product[47]) );
  OAI22X1TS U1028 ( .A0(n821), .A1(n1020), .B0(n80), .B1(n807), .Y(n811) );
  OAI22X1TS U1029 ( .A0(n808), .A1(n882), .B0(n820), .B1(n884), .Y(n810) );
  OAI21XLTS U1030 ( .A0(n811), .A1(n810), .B0(n76), .Y(n809) );
  OAI31X1TS U1031 ( .A0(n811), .A1(n76), .A2(n810), .B0(n809), .Y(
        \mult_x_1/n1216 ) );
  OAI22X1TS U1032 ( .A0(n819), .A1(n1020), .B0(n80), .B1(n812), .Y(n815) );
  OAI22X1TS U1033 ( .A0(n821), .A1(n818), .B0(n820), .B1(n882), .Y(n814) );
  OAI21XLTS U1034 ( .A0(n815), .A1(n814), .B0(n76), .Y(n813) );
  OAI31X1TS U1035 ( .A0(n815), .A1(n76), .A2(n814), .B0(n813), .Y(
        \mult_x_1/n1217 ) );
  OAI22X1TS U1036 ( .A0(n817), .A1(n1020), .B0(n816), .B1(n80), .Y(n824) );
  OAI22X1TS U1037 ( .A0(n821), .A1(n820), .B0(n819), .B1(n818), .Y(n823) );
  OAI21XLTS U1038 ( .A0(n824), .A1(n823), .B0(n76), .Y(n822) );
  OAI31X1TS U1039 ( .A0(n824), .A1(n76), .A2(n823), .B0(n822), .Y(
        \mult_x_1/n1218 ) );
  INVX2TS U1040 ( .A(n828), .Y(Product[48]) );
  OAI22X1TS U1041 ( .A0(n1023), .A1(n1009), .B0(n93), .B1(n1001), .Y(n830) );
  OAI21XLTS U1042 ( .A0(n970), .A1(n830), .B0(n1028), .Y(n829) );
  OAI31X1TS U1043 ( .A0(n970), .A1(n1028), .A2(n830), .B0(n829), .Y(
        \mult_x_1/n1232 ) );
  OAI22X1TS U1044 ( .A0(n1023), .A1(n831), .B0(n93), .B1(n992), .Y(n834) );
  OAI22X1TS U1045 ( .A0(n906), .A1(n996), .B0(n904), .B1(\mult_x_1/n404 ), .Y(
        n833) );
  OAI21XLTS U1046 ( .A0(n834), .A1(n833), .B0(n1028), .Y(n832) );
  OAI31X1TS U1047 ( .A0(n834), .A1(n1028), .A2(n833), .B0(n832), .Y(
        \mult_x_1/n1235 ) );
  OAI22X1TS U1048 ( .A0(n1023), .A1(n835), .B0(n93), .B1(\mult_x_1/n404 ), .Y(
        n838) );
  OAI22X1TS U1049 ( .A0(n906), .A1(n1001), .B0(n904), .B1(n996), .Y(n837) );
  OAI21XLTS U1050 ( .A0(n838), .A1(n837), .B0(n1028), .Y(n836) );
  OAI31X1TS U1051 ( .A0(n838), .A1(n1028), .A2(n837), .B0(n836), .Y(
        \mult_x_1/n1234 ) );
  OAI22X1TS U1052 ( .A0(n1023), .A1(n839), .B0(n93), .B1(n895), .Y(n842) );
  OAI22X1TS U1053 ( .A0(n906), .A1(n1030), .B0(n904), .B1(n896), .Y(n841) );
  OAI21XLTS U1054 ( .A0(n842), .A1(n841), .B0(n1028), .Y(n840) );
  OAI31X1TS U1055 ( .A0(n842), .A1(n1028), .A2(n841), .B0(n840), .Y(
        \mult_x_1/n1243 ) );
  OAI22X1TS U1056 ( .A0(n1023), .A1(n843), .B0(n93), .B1(n852), .Y(n846) );
  OAI22X1TS U1057 ( .A0(n906), .A1(n877), .B0(n904), .B1(n864), .Y(n845) );
  OAI21XLTS U1058 ( .A0(n846), .A1(n845), .B0(n1028), .Y(n844) );
  OAI31X1TS U1059 ( .A0(n846), .A1(n1028), .A2(n845), .B0(n844), .Y(
        \mult_x_1/n1247 ) );
  OAI22X1TS U1060 ( .A0(n1023), .A1(n847), .B0(n93), .B1(n885), .Y(n850) );
  OAI22X1TS U1061 ( .A0(n906), .A1(n864), .B0(n904), .B1(n852), .Y(n849) );
  OAI21XLTS U1062 ( .A0(n850), .A1(n849), .B0(n1028), .Y(n848) );
  OAI31X1TS U1063 ( .A0(n850), .A1(n1028), .A2(n849), .B0(n848), .Y(
        \mult_x_1/n1248 ) );
  OAI22X1TS U1064 ( .A0(n1023), .A1(n851), .B0(n93), .B1(n884), .Y(n855) );
  OAI22X1TS U1065 ( .A0(n906), .A1(n852), .B0(n904), .B1(n885), .Y(n854) );
  OAI21XLTS U1066 ( .A0(n855), .A1(n854), .B0(n1028), .Y(n853) );
  OAI31X1TS U1067 ( .A0(n855), .A1(n1028), .A2(n854), .B0(n853), .Y(
        \mult_x_1/n1249 ) );
  OAI22X1TS U1068 ( .A0(n1023), .A1(n856), .B0(n93), .B1(n905), .Y(n859) );
  OAI22X1TS U1069 ( .A0(n906), .A1(n992), .B0(n904), .B1(n988), .Y(n858) );
  OAI21XLTS U1070 ( .A0(n859), .A1(n858), .B0(n1028), .Y(n857) );
  OAI31X1TS U1071 ( .A0(n859), .A1(n1028), .A2(n858), .B0(n857), .Y(
        \mult_x_1/n1237 ) );
  OAI22X1TS U1072 ( .A0(n1023), .A1(n860), .B0(n93), .B1(n1030), .Y(n863) );
  OAI22X1TS U1073 ( .A0(n906), .A1(n977), .B0(n904), .B1(n973), .Y(n862) );
  OAI21XLTS U1074 ( .A0(n863), .A1(n862), .B0(n1028), .Y(n861) );
  OAI31X1TS U1075 ( .A0(n863), .A1(n1028), .A2(n862), .B0(n861), .Y(
        \mult_x_1/n1241 ) );
  OAI22X1TS U1076 ( .A0(n1023), .A1(n865), .B0(n93), .B1(n864), .Y(n868) );
  OAI22X1TS U1077 ( .A0(n906), .A1(n893), .B0(n904), .B1(n877), .Y(n867) );
  OAI21XLTS U1078 ( .A0(n868), .A1(n867), .B0(n1028), .Y(n866) );
  OAI31X1TS U1079 ( .A0(n868), .A1(n1028), .A2(n867), .B0(n866), .Y(
        \mult_x_1/n1246 ) );
  OAI22X1TS U1080 ( .A0(n1023), .A1(n869), .B0(n93), .B1(n903), .Y(n872) );
  OAI22X1TS U1081 ( .A0(n906), .A1(n988), .B0(n904), .B1(n905), .Y(n871) );
  OAI21XLTS U1082 ( .A0(n872), .A1(n871), .B0(n1028), .Y(n870) );
  OAI31X1TS U1083 ( .A0(n872), .A1(n1028), .A2(n871), .B0(n870), .Y(
        \mult_x_1/n1238 ) );
  OAI22X1TS U1084 ( .A0(n1023), .A1(n873), .B0(n93), .B1(n896), .Y(n876) );
  OAI22X1TS U1085 ( .A0(n906), .A1(n973), .B0(n904), .B1(n1030), .Y(n875) );
  OAI21XLTS U1086 ( .A0(n876), .A1(n875), .B0(n1028), .Y(n874) );
  OAI31X1TS U1087 ( .A0(n876), .A1(n1028), .A2(n875), .B0(n874), .Y(
        \mult_x_1/n1242 ) );
  OAI22X1TS U1088 ( .A0(n1023), .A1(n878), .B0(n93), .B1(n877), .Y(n881) );
  OAI22X1TS U1089 ( .A0(n906), .A1(n895), .B0(n904), .B1(n893), .Y(n880) );
  OAI21XLTS U1090 ( .A0(n881), .A1(n880), .B0(n1028), .Y(n879) );
  OAI31X1TS U1091 ( .A0(n881), .A1(n1028), .A2(n880), .B0(n879), .Y(
        \mult_x_1/n1245 ) );
  OAI22X1TS U1092 ( .A0(n1023), .A1(n883), .B0(n93), .B1(n882), .Y(n888) );
  OAI22X1TS U1093 ( .A0(n906), .A1(n885), .B0(n904), .B1(n884), .Y(n887) );
  OAI21XLTS U1094 ( .A0(n888), .A1(n887), .B0(n1028), .Y(n886) );
  OAI31X1TS U1095 ( .A0(n888), .A1(n1028), .A2(n887), .B0(n886), .Y(
        \mult_x_1/n1250 ) );
  OAI22X1TS U1096 ( .A0(n1023), .A1(n889), .B0(n93), .B1(n988), .Y(n892) );
  OAI22X1TS U1097 ( .A0(n906), .A1(\mult_x_1/n404 ), .B0(n904), .B1(n992), .Y(
        n891) );
  OAI21XLTS U1098 ( .A0(n892), .A1(n891), .B0(n1028), .Y(n890) );
  OAI31X1TS U1099 ( .A0(n892), .A1(n1028), .A2(n891), .B0(n890), .Y(
        \mult_x_1/n1236 ) );
  OAI22X1TS U1100 ( .A0(n1023), .A1(n894), .B0(n93), .B1(n893), .Y(n899) );
  OAI22X1TS U1101 ( .A0(n906), .A1(n896), .B0(n904), .B1(n895), .Y(n898) );
  OAI21XLTS U1102 ( .A0(n899), .A1(n898), .B0(n1028), .Y(n897) );
  OAI31X1TS U1103 ( .A0(n899), .A1(n1028), .A2(n898), .B0(n897), .Y(
        \mult_x_1/n1244 ) );
  OAI22X1TS U1104 ( .A0(n1023), .A1(n981), .B0(n93), .B1(n973), .Y(n902) );
  OAI22X1TS U1105 ( .A0(n906), .A1(n903), .B0(n904), .B1(n977), .Y(n901) );
  OAI21XLTS U1106 ( .A0(n902), .A1(n901), .B0(n1028), .Y(n900) );
  OAI31X1TS U1107 ( .A0(n902), .A1(n1028), .A2(n901), .B0(n900), .Y(
        \mult_x_1/n1240 ) );
  OAI22X1TS U1108 ( .A0(n1023), .A1(n985), .B0(n93), .B1(n977), .Y(n909) );
  OAI22X1TS U1109 ( .A0(n906), .A1(n905), .B0(n904), .B1(n903), .Y(n908) );
  OAI21XLTS U1110 ( .A0(n909), .A1(n908), .B0(n1028), .Y(n907) );
  OAI31X1TS U1111 ( .A0(n909), .A1(n1028), .A2(n908), .B0(n907), .Y(
        \mult_x_1/n1239 ) );
  INVX2TS U1112 ( .A(n913), .Y(\mult_x_1/n796 ) );
  INVX2TS U1113 ( .A(n914), .Y(Product[63]) );
  OA21XLTS U1114 ( .A0(n924), .A1(n923), .B0(n922), .Y(Product[3]) );
  NAND2X1TS U1115 ( .A(A[2]), .B(Product[0]), .Y(n926) );
  OA21XLTS U1116 ( .A0(n927), .A1(n926), .B0(n925), .Y(Product[1]) );
  AOI2BB2XLTS U1117 ( .B0(n929), .B1(n928), .A0N(n928), .A1N(n929), .Y(n930)
         );
  XNOR2X1TS U1118 ( .A(n931), .B(n930), .Y(\mult_x_1/n670 ) );
  AOI21X1TS U1119 ( .A0(n933), .A1(n932), .B0(n931), .Y(\mult_x_1/n683 ) );
  OA21XLTS U1120 ( .A0(n935), .A1(n934), .B0(n933), .Y(\mult_x_1/n694 ) );
  OAI31X1TS U1121 ( .A0(n937), .A1(n939), .A2(n1016), .B0(n936), .Y(n938) );
  AOI21X1TS U1122 ( .A0(n939), .A1(n1016), .B0(n938), .Y(\mult_x_1/n743 ) );
  OAI31X1TS U1123 ( .A0(n941), .A1(n943), .A2(n957), .B0(n940), .Y(n942) );
  AOI21X1TS U1124 ( .A0(n943), .A1(n957), .B0(n942), .Y(\mult_x_1/n785 ) );
  OAI22X1TS U1125 ( .A0(n967), .A1(n1012), .B0(n1011), .B1(n996), .Y(n944) );
  AOI211XLTS U1126 ( .A0(n946), .A1(B[22]), .B0(n945), .C0(n944), .Y(n947) );
  XNOR2X1TS U1127 ( .A(A[20]), .B(n947), .Y(\mult_x_1/n1058 ) );
  OAI22X1TS U1128 ( .A0(n967), .A1(n404), .B0(n1014), .B1(n996), .Y(n948) );
  AOI211XLTS U1129 ( .A0(n950), .A1(B[22]), .B0(n949), .C0(n948), .Y(n951) );
  XNOR2X1TS U1130 ( .A(A[17]), .B(n951), .Y(\mult_x_1/n1093 ) );
  OAI22X1TS U1131 ( .A0(n967), .A1(n1018), .B0(n1017), .B1(n996), .Y(n952) );
  AOI211XLTS U1132 ( .A0(n954), .A1(B[22]), .B0(n953), .C0(n952), .Y(n955) );
  XNOR2X1TS U1133 ( .A(A[14]), .B(n955), .Y(\mult_x_1/n1128 ) );
  OAI21XLTS U1134 ( .A0(n652), .A1(n1022), .B0(n958), .Y(n956) );
  XNOR2X1TS U1135 ( .A(n957), .B(n956), .Y(\mult_x_1/n1161 ) );
  OAI22X1TS U1136 ( .A0(n967), .A1(n652), .B0(n958), .B1(n996), .Y(n959) );
  AOI211XLTS U1137 ( .A0(n961), .A1(B[22]), .B0(n960), .C0(n959), .Y(n962) );
  XNOR2X1TS U1138 ( .A(A[11]), .B(n962), .Y(\mult_x_1/n1163 ) );
  OAI22X1TS U1139 ( .A0(n967), .A1(n80), .B0(n1020), .B1(n996), .Y(n963) );
  AOI211XLTS U1140 ( .A0(n965), .A1(B[22]), .B0(n964), .C0(n963), .Y(n966) );
  XNOR2X1TS U1141 ( .A(A[8]), .B(n966), .Y(\mult_x_1/n1198 ) );
  OAI22X1TS U1142 ( .A0(n967), .A1(n1023), .B0(n93), .B1(n996), .Y(n968) );
  AOI211XLTS U1143 ( .A0(n970), .A1(B[22]), .B0(n969), .C0(n968), .Y(n971) );
  XNOR2X1TS U1144 ( .A(n1036), .B(n971), .Y(\mult_x_1/n1233 ) );
  AOI22X1TS U1145 ( .A0(n1008), .A1(B[12]), .B0(n999), .B1(B[13]), .Y(n972) );
  OAI21XLTS U1146 ( .A0(n1002), .A1(n973), .B0(n972), .Y(n974) );
  AOI21X1TS U1147 ( .A0(n1010), .A1(n975), .B0(n974), .Y(\mult_x_1/n1032 ) );
  AOI22X1TS U1148 ( .A0(n1008), .A1(B[13]), .B0(n999), .B1(B[14]), .Y(n976) );
  OAI21XLTS U1149 ( .A0(n1002), .A1(n977), .B0(n976), .Y(n978) );
  AOI21X1TS U1150 ( .A0(n1010), .A1(n979), .B0(n978), .Y(\mult_x_1/n1031 ) );
  AOI22X1TS U1151 ( .A0(n983), .A1(B[16]), .B0(n1008), .B1(B[14]), .Y(n980) );
  OAI21XLTS U1152 ( .A0(n1006), .A1(n981), .B0(n980), .Y(n982) );
  AOI21X1TS U1153 ( .A0(n999), .A1(B[15]), .B0(n982), .Y(\mult_x_1/n1030 ) );
  AOI22X1TS U1154 ( .A0(n983), .A1(B[17]), .B0(n999), .B1(B[16]), .Y(n984) );
  OAI21XLTS U1155 ( .A0(n1006), .A1(n985), .B0(n984), .Y(n986) );
  AOI21X1TS U1156 ( .A0(n1008), .A1(B[15]), .B0(n986), .Y(\mult_x_1/n1029 ) );
  AOI22X1TS U1157 ( .A0(n1008), .A1(B[16]), .B0(n999), .B1(B[17]), .Y(n987) );
  OAI21XLTS U1158 ( .A0(n1002), .A1(n988), .B0(n987), .Y(n989) );
  AOI21X1TS U1159 ( .A0(n1010), .A1(n990), .B0(n989), .Y(\mult_x_1/n1028 ) );
  AOI22X1TS U1160 ( .A0(n1008), .A1(B[17]), .B0(n999), .B1(B[18]), .Y(n991) );
  OAI21XLTS U1161 ( .A0(n1002), .A1(n992), .B0(n991), .Y(n993) );
  AOI21X1TS U1162 ( .A0(n1010), .A1(n994), .B0(n993), .Y(\mult_x_1/n1027 ) );
  AOI22X1TS U1163 ( .A0(n1008), .A1(B[19]), .B0(n999), .B1(B[20]), .Y(n995) );
  OAI21XLTS U1164 ( .A0(n1002), .A1(n996), .B0(n995), .Y(n997) );
  AOI21X1TS U1165 ( .A0(n1010), .A1(n998), .B0(n997), .Y(\mult_x_1/n1025 ) );
  AOI22X1TS U1166 ( .A0(n1008), .A1(B[20]), .B0(n999), .B1(B[21]), .Y(n1000)
         );
  OAI21XLTS U1167 ( .A0(n1002), .A1(n1001), .B0(n1000), .Y(n1003) );
  AOI21X1TS U1168 ( .A0(n1010), .A1(n1004), .B0(n1003), .Y(\mult_x_1/n1024 )
         );
  OAI21XLTS U1169 ( .A0(n1006), .A1(n1009), .B0(n1005), .Y(n1007) );
  AOI21X1TS U1170 ( .A0(n1008), .A1(B[22]), .B0(n1007), .Y(\mult_x_1/n1022 )
         );
  AOI21X1TS U1171 ( .A0(n1010), .A1(n1009), .B0(n1008), .Y(\mult_x_1/n1021 )
         );
  OAI21XLTS U1172 ( .A0(n1012), .A1(n1022), .B0(n1011), .Y(n1013) );
  XNOR2X1TS U1173 ( .A(n917), .B(n1013), .Y(\mult_x_1/n1056 ) );
  OAI21XLTS U1174 ( .A0(n404), .A1(n1022), .B0(n1014), .Y(n1015) );
  XNOR2X1TS U1175 ( .A(n1016), .B(n1015), .Y(\mult_x_1/n1091 ) );
  OAI21XLTS U1176 ( .A0(n1018), .A1(n1022), .B0(n1017), .Y(n1019) );
  XNOR2X1TS U1177 ( .A(n1035), .B(n1019), .Y(\mult_x_1/n1126 ) );
  OAI21XLTS U1178 ( .A0(n80), .A1(n1022), .B0(n1020), .Y(n1021) );
  XNOR2X1TS U1179 ( .A(n76), .B(n1021), .Y(\mult_x_1/n1196 ) );
  OAI21XLTS U1180 ( .A0(n1023), .A1(n1022), .B0(n93), .Y(n1024) );
  XNOR2X1TS U1181 ( .A(n1028), .B(n1024), .Y(\mult_x_1/n1231 ) );
  AOI21X1TS U1182 ( .A0(A[8]), .A1(n1026), .B0(n1025), .Y(\mult_x_1/n452 ) );
  OAI21XLTS U1183 ( .A0(n1028), .A1(n1027), .B0(n1026), .Y(n1029) );
  AOI21X1TS U1184 ( .A0(n1030), .A1(n1029), .B0(\mult_x_1/n463 ), .Y(
        \mult_x_1/n491 ) );
endmodule


module mux2_1_1 ( selector, data_in_0, data_in_1, data_out );
  input [31:0] data_in_0;
  input [31:0] data_in_1;
  output [31:0] data_out;
  input selector;
  wire   n1, n2;

  INVX2TS U1 ( .A(selector), .Y(n1) );
  INVX2TS U2 ( .A(n1), .Y(n2) );
  AO22XLTS U3 ( .A0(n2), .A1(data_in_1[11]), .B0(n1), .B1(data_in_0[11]), .Y(
        data_out[11]) );
  AO22XLTS U4 ( .A0(n2), .A1(data_in_1[5]), .B0(n1), .B1(data_in_0[5]), .Y(
        data_out[5]) );
  AO22XLTS U5 ( .A0(n2), .A1(data_in_1[17]), .B0(n1), .B1(data_in_0[17]), .Y(
        data_out[17]) );
  AO22XLTS U6 ( .A0(n2), .A1(data_in_1[23]), .B0(n1), .B1(data_in_0[23]), .Y(
        data_out[23]) );
  AO22XLTS U7 ( .A0(n2), .A1(data_in_1[8]), .B0(n1), .B1(data_in_0[8]), .Y(
        data_out[8]) );
  AO22XLTS U8 ( .A0(n2), .A1(data_in_1[14]), .B0(n1), .B1(data_in_0[14]), .Y(
        data_out[14]) );
  AO22XLTS U9 ( .A0(n2), .A1(data_in_1[20]), .B0(n1), .B1(data_in_0[20]), .Y(
        data_out[20]) );
  AO22XLTS U10 ( .A0(n2), .A1(data_in_1[26]), .B0(n1), .B1(data_in_0[26]), .Y(
        data_out[26]) );
  AO22XLTS U11 ( .A0(n2), .A1(data_in_1[29]), .B0(n1), .B1(data_in_0[29]), .Y(
        data_out[29]) );
  AO22XLTS U12 ( .A0(n2), .A1(data_in_1[0]), .B0(n1), .B1(data_in_0[0]), .Y(
        data_out[0]) );
  AO22XLTS U13 ( .A0(n2), .A1(data_in_1[1]), .B0(n1), .B1(data_in_0[1]), .Y(
        data_out[1]) );
  AO22XLTS U14 ( .A0(n2), .A1(data_in_1[3]), .B0(n1), .B1(data_in_0[3]), .Y(
        data_out[3]) );
  AO22XLTS U15 ( .A0(n2), .A1(data_in_1[4]), .B0(n1), .B1(data_in_0[4]), .Y(
        data_out[4]) );
  AO22XLTS U16 ( .A0(n2), .A1(data_in_1[6]), .B0(n1), .B1(data_in_0[6]), .Y(
        data_out[6]) );
  AO22XLTS U17 ( .A0(n2), .A1(data_in_1[7]), .B0(n1), .B1(data_in_0[7]), .Y(
        data_out[7]) );
  AO22XLTS U18 ( .A0(n2), .A1(data_in_1[30]), .B0(n1), .B1(data_in_0[30]), .Y(
        data_out[30]) );
  AO22XLTS U19 ( .A0(n2), .A1(data_in_1[2]), .B0(n1), .B1(data_in_0[2]), .Y(
        data_out[2]) );
  AO22XLTS U20 ( .A0(n2), .A1(data_in_1[9]), .B0(n1), .B1(data_in_0[9]), .Y(
        data_out[9]) );
  AO22XLTS U21 ( .A0(n2), .A1(data_in_1[10]), .B0(n1), .B1(data_in_0[10]), .Y(
        data_out[10]) );
  AO22XLTS U22 ( .A0(n2), .A1(data_in_1[12]), .B0(n1), .B1(data_in_0[12]), .Y(
        data_out[12]) );
  AO22XLTS U23 ( .A0(n2), .A1(data_in_1[13]), .B0(n1), .B1(data_in_0[13]), .Y(
        data_out[13]) );
  AO22XLTS U24 ( .A0(n2), .A1(data_in_1[15]), .B0(n1), .B1(data_in_0[15]), .Y(
        data_out[15]) );
  AO22XLTS U25 ( .A0(n2), .A1(data_in_1[16]), .B0(n1), .B1(data_in_0[16]), .Y(
        data_out[16]) );
  AO22XLTS U26 ( .A0(n2), .A1(data_in_1[18]), .B0(n1), .B1(data_in_0[18]), .Y(
        data_out[18]) );
  AO22XLTS U27 ( .A0(n2), .A1(data_in_1[19]), .B0(n1), .B1(data_in_0[19]), .Y(
        data_out[19]) );
  AO22XLTS U28 ( .A0(n2), .A1(data_in_1[21]), .B0(n1), .B1(data_in_0[21]), .Y(
        data_out[21]) );
  AO22XLTS U29 ( .A0(n2), .A1(data_in_1[22]), .B0(n1), .B1(data_in_0[22]), .Y(
        data_out[22]) );
  AO22XLTS U30 ( .A0(n2), .A1(data_in_1[24]), .B0(n1), .B1(data_in_0[24]), .Y(
        data_out[24]) );
  AO22XLTS U31 ( .A0(n2), .A1(data_in_1[25]), .B0(n1), .B1(data_in_0[25]), .Y(
        data_out[25]) );
  AO22XLTS U32 ( .A0(n2), .A1(data_in_1[31]), .B0(n1), .B1(data_in_0[31]), .Y(
        data_out[31]) );
  AO22XLTS U33 ( .A0(n2), .A1(data_in_1[27]), .B0(n1), .B1(data_in_0[27]), .Y(
        data_out[27]) );
  AO22XLTS U34 ( .A0(n2), .A1(data_in_1[28]), .B0(n1), .B1(data_in_0[28]), .Y(
        data_out[28]) );
endmodule


module calculator ( clk, start, reset, mode, calculator_input, n_input, 
        regacc_out, state_out, Coutadd, Coutone, Couttwo, m14_out, alutwo_out, 
        m17_out, m18_out, srmq_out, regec_out, regeb_out, rf_aout, regi_out, 
        regcurrterm_out, regsum_out, srmt_out, regms_out, reges_out, reget_out, 
        regss0_out, reges0_out, ssrms0_out, aluone_out, regreg_out, rege_out
 );
  input [2:0] mode;
  input [31:0] calculator_input;
  input [31:0] n_input;
  output [31:0] regacc_out;
  output [8:0] state_out;
  output [31:0] m14_out;
  output [31:0] alutwo_out;
  output [31:0] m17_out;
  output [31:0] m18_out;
  output [63:0] srmq_out;
  output [31:0] regec_out;
  output [31:0] regeb_out;
  output [31:0] rf_aout;
  output [5:0] regi_out;
  output [31:0] regcurrterm_out;
  output [31:0] regsum_out;
  output [31:0] srmt_out;
  output [31:0] regms_out;
  output [31:0] reges_out;
  output [31:0] reget_out;
  output [31:0] reges0_out;
  output [63:0] ssrms0_out;
  output [31:0] aluone_out;
  output [31:0] regreg_out;
  output [31:0] rege_out;
  input clk, start, reset;
  output Coutadd, Coutone, Couttwo, regss0_out;
  wire   n4821, regsp_out, mux5, \m6_out[0] , regst_out, mux7, mux10, mux11,
         mux15, regsc_out, regsa_out, mux19, \mux20[0] , mux22, mux23,
         regsq_out, reg_ss, regss_out, reg_st, reg_ss0, reg_sc, reg_sb,
         regsb_out, reg_sa, reg_sp, reg_i, reg_index, reg_es, reg_et, reg_acc,
         reg_sum, reg_currterm, reg_numbit, reg_es0, reg_e, reg_ec, reg_eb,
         reg_mb, reg_ea, reg_ma, \sr_mt[0] , sumorrr_out, xor3_out, rf_reb,
         rf_rea, \comp1/N0 , \comp2/N0 , \aluone/N325 , \aluone/N324 ,
         \alutwo/N325 , \alutwo/N324 , \count/N34 , \count/N32 , \count/N30 ,
         \count/N29 , \C43/DATA3_1 , \C43/DATA3_2 , \C43/DATA3_3 ,
         \C43/DATA3_4 , n1649, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, \DP_OP_117J3_124_765/n2 ,
         \DP_OP_117J3_124_765/n3 , \DP_OP_117J3_124_765/n4 ,
         \DP_OP_117J3_124_765/n5 , n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4819;
  wire   [31:0] m1_out;
  wire   [2:0] mux2;
  wire   [31:0] m2_out;
  wire   [2:0] mux3;
  wire   [31:0] m3_out;
  wire   [63:0] srmp_out;
  wire   [1:0] mux4;
  wire   [31:0] bs2_out;
  wire   [31:0] regr_out;
  wire   [31:0] m4_out;
  wire   [31:0] m5_out;
  wire   [1:0] mux6;
  wire   [2:0] mux8;
  wire   [2:0] mux9;
  wire   [31:0] m10_out;
  wire   [1:0] mux12;
  wire   [63:0] mult1_out;
  wire   [2:0] mux13;
  wire   [5:0] m13_out;
  wire   [1:0] mux14;
  wire   [5:0] rf_rab;
  wire   [5:0] regindex_out;
  wire   [5:0] m15_out;
  wire   [2:0] mux17;
  wire   [31:0] regeq_out;
  wire   [31:0] regep_out;
  wire   [31:0] regea_out;
  wire   [31:0] regma_out;
  wire   [31:0] regmc_out;
  wire   [31:0] m19_out;
  wire   [31:0] regres_out;
  wire   [1:0] mux21;
  wire   [31:0] rf_bout;
  wire   [31:0] regnumbit_out;
  wire   [5:0] pe_out;
  wire   [31:0] regmb_out;
  wire   [1:0] sr_res;
  wire   [1:0] sr_mp;
  wire   [63:0] mult2_out;
  wire   [1:0] sr_mq;
  wire   [2:0] ssr_ms0;
  wire   [5:0] count_out;
  wire   [2:0] alu1;
  wire   [2:0] alu2;
  wire   [2:0] counterii;
  wire   [5:0] rf_wa;
  wire   [5:0] rf_raa;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25;

  mux4_1_0 m4 ( .selector(mux4), .data_in_00(bs2_out), .data_in_01(regr_out), 
        .data_in_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        regsum_out[22:0]}), .data_in_11({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .data_out(m4_out) );
  mux2_1_0 m5 ( .selector(mux5), .data_in_0(bs2_out), .data_in_1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, regcurrterm_out[22:0]}), 
        .data_out(m5_out) );
  mux2_1_1 m10 ( .selector(mux10), .data_in_0(srmt_out), .data_in_1(regms_out), 
        .data_out(m10_out) );
  register_0 regnumbit ( .clk(clk), .load(reg_numbit), .data_in(aluone_out), 
        .data_out(regnumbit_out) );
  mult32_0 mult1 ( .A(regms_out), .B(srmt_out), .Product(mult1_out) );
  mult32_1 mult2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        regmb_out[22:18], n4816, regmb_out[16:12], n4815, regmb_out[10:3], 
        n4814, regmb_out[1:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1, m19_out[22:0]}), .Product({mult2_out[63], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, mult2_out[53:0]}) );
  Bshifterright bs2 ( .data_in(m10_out), .data_out(bs2_out), .bits(
        regnumbit_out) );
  RF rf ( .clk(clk), .data_in(m14_out), .data_outA(rf_aout), .data_outB(
        rf_bout), .WA({rf_wa[5], 1'b0, 1'b0, 1'b0, rf_wa[1:0]}), .RAA({
        rf_raa[5], 1'b0, 1'b0, 1'b0, rf_raa[1:0]}), .RAB(m15_out), .enable({
        1'b0, rf_reb, rf_rea}) );
  FSM FSM ( .clk(clk), .reset(reset), .start(start), .mq47(srmq_out[47]), 
        .mp47(srmp_out[47]), .r31(regr_out[31]), .msb(count_out[5]), .ms0_24(
        ssrms0_out[24]), .ms0_23(ssrms0_out[23]), .ms0_63(ssrms0_out[63]), 
        .comp1_g(\comp1/N0 ), .comp2_g(\comp2/N0 ), .stxor(xor3_out), .st(
        regst_out), .sumor(sumorrr_out), .mode(mode), .mux5(mux5), .mux7(mux7), 
        .mux10(mux10), .mux11(mux11), .mux15(mux15), .mux19(mux19), .mux22(
        mux22), .mux23(mux23), .mux1({SYNOPSYS_UNCONNECTED__9, n1992}), .mux4(
        mux4), .mux6(mux6), .mux12(mux12), .mux14({n1991, mux14[0]}), .mux20({
        SYNOPSYS_UNCONNECTED__10, \mux20[0] }), .mux21(mux21), .mux2(mux2), 
        .mux3({mux3[2:1], SYNOPSYS_UNCONNECTED__11}), .mux8({mux8[2], 
        SYNOPSYS_UNCONNECTED__12, mux8[0]}), .mux9(mux9), .mux13(mux13), 
        .mux17({mux17[2], SYNOPSYS_UNCONNECTED__13, mux17[0]}), .rf_rea(rf_rea), .rf_reb(rf_reb), .rf_wa({rf_wa[5], SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, rf_wa[1:0]}), 
        .rf_raa({rf_raa[5], SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, rf_raa[1:0]}), .rf_rab({rf_rab[5], 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, rf_rab[1:0]}), .reg_sum(reg_sum), .reg_i(
        reg_i), .reg_currterm(reg_currterm), .reg_index(reg_index), .reg_reg(
        n1994), .reg_r(n1993), .reg_numbit(reg_numbit), .reg_e(reg_e), 
        .reg_acc(reg_acc), .reg_sc(reg_sc), .reg_ec(reg_ec), .reg_mc(n1990), 
        .reg_sb(reg_sb), .reg_eb(reg_eb), .reg_mb(reg_mb), .reg_sa(reg_sa), 
        .reg_ea(reg_ea), .reg_ma(reg_ma), .reg_eq(n1988), .reg_ss(reg_ss), 
        .reg_es(reg_es), .reg_ms(n1989), .reg_st(reg_st), .reg_et(reg_et), 
        .reg_sp(reg_sp), .reg_ep(n1986), .reg_es0(reg_es0), .reg_ss0(reg_ss0), 
        .sr_res(sr_res), .sr_mq(sr_mq), .sr_mt({SYNOPSYS_UNCONNECTED__23, 
        \sr_mt[0] }), .sr_mp(sr_mp), .ssr_ms0({SYNOPSYS_UNCONNECTED__24, 
        ssr_ms0[1:0]}), .alu1({\aluone/N324 , alu1[1:0]}), .alu2({
        \alutwo/N324 , alu2[1:0]}), .counterii({counterii[2:1], 
        SYNOPSYS_UNCONNECTED__25}), .state(state_out) );
  EDFFX1TS \regep/data_out_buffer_reg[0]  ( .D(alutwo_out[0]), .E(n1986), .CK(
        clk), .Q(regep_out[0]) );
  EDFFX1TS \regep/data_out_buffer_reg[1]  ( .D(alutwo_out[1]), .E(n1986), .CK(
        clk), .Q(regep_out[1]) );
  EDFFX1TS \regep/data_out_buffer_reg[2]  ( .D(alutwo_out[2]), .E(n1986), .CK(
        clk), .Q(regep_out[2]) );
  EDFFX1TS \regep/data_out_buffer_reg[3]  ( .D(alutwo_out[3]), .E(n1986), .CK(
        clk), .Q(regep_out[3]) );
  EDFFX1TS \regep/data_out_buffer_reg[4]  ( .D(alutwo_out[4]), .E(n1986), .CK(
        clk), .Q(regep_out[4]) );
  EDFFX1TS \regep/data_out_buffer_reg[5]  ( .D(alutwo_out[5]), .E(n1986), .CK(
        clk), .Q(regep_out[5]) );
  EDFFX1TS \regep/data_out_buffer_reg[6]  ( .D(alutwo_out[6]), .E(n1986), .CK(
        clk), .Q(regep_out[6]) );
  EDFFX1TS \regep/data_out_buffer_reg[7]  ( .D(alutwo_out[7]), .E(n1986), .CK(
        clk), .Q(regep_out[7]) );
  EDFFX1TS \regep/data_out_buffer_reg[8]  ( .D(alutwo_out[8]), .E(n1986), .CK(
        clk), .Q(regep_out[8]) );
  EDFFX1TS \regep/data_out_buffer_reg[9]  ( .D(alutwo_out[9]), .E(n1986), .CK(
        clk), .Q(regep_out[9]) );
  EDFFX1TS \regep/data_out_buffer_reg[10]  ( .D(alutwo_out[10]), .E(n1986), 
        .CK(clk), .Q(regep_out[10]) );
  EDFFX1TS \regep/data_out_buffer_reg[11]  ( .D(alutwo_out[11]), .E(n1986), 
        .CK(clk), .Q(regep_out[11]) );
  EDFFX1TS \regep/data_out_buffer_reg[12]  ( .D(alutwo_out[12]), .E(n1986), 
        .CK(clk), .Q(regep_out[12]) );
  EDFFX1TS \regep/data_out_buffer_reg[13]  ( .D(alutwo_out[13]), .E(n1986), 
        .CK(clk), .Q(regep_out[13]) );
  EDFFX1TS \regep/data_out_buffer_reg[14]  ( .D(alutwo_out[14]), .E(n1986), 
        .CK(clk), .Q(regep_out[14]) );
  EDFFX1TS \regep/data_out_buffer_reg[15]  ( .D(alutwo_out[15]), .E(n1986), 
        .CK(clk), .Q(regep_out[15]) );
  EDFFX1TS \regep/data_out_buffer_reg[16]  ( .D(alutwo_out[16]), .E(n1986), 
        .CK(clk), .Q(regep_out[16]) );
  EDFFX1TS \regep/data_out_buffer_reg[17]  ( .D(alutwo_out[17]), .E(n1986), 
        .CK(clk), .Q(regep_out[17]) );
  EDFFX1TS \regep/data_out_buffer_reg[18]  ( .D(alutwo_out[18]), .E(n1986), 
        .CK(clk), .Q(regep_out[18]) );
  EDFFX1TS \regep/data_out_buffer_reg[19]  ( .D(alutwo_out[19]), .E(n1986), 
        .CK(clk), .Q(regep_out[19]) );
  EDFFX1TS \regep/data_out_buffer_reg[20]  ( .D(alutwo_out[20]), .E(n1986), 
        .CK(clk), .Q(regep_out[20]) );
  EDFFX1TS \regep/data_out_buffer_reg[21]  ( .D(alutwo_out[21]), .E(n1986), 
        .CK(clk), .Q(regep_out[21]) );
  EDFFX1TS \regep/data_out_buffer_reg[22]  ( .D(alutwo_out[22]), .E(n1986), 
        .CK(clk), .Q(regep_out[22]) );
  EDFFX1TS \regep/data_out_buffer_reg[23]  ( .D(alutwo_out[23]), .E(n1986), 
        .CK(clk), .Q(regep_out[23]) );
  EDFFX1TS \regep/data_out_buffer_reg[24]  ( .D(alutwo_out[24]), .E(n1986), 
        .CK(clk), .Q(regep_out[24]) );
  EDFFX1TS \regep/data_out_buffer_reg[25]  ( .D(alutwo_out[25]), .E(n1986), 
        .CK(clk), .Q(regep_out[25]) );
  EDFFX1TS \regep/data_out_buffer_reg[26]  ( .D(alutwo_out[26]), .E(n1986), 
        .CK(clk), .Q(regep_out[26]) );
  EDFFX1TS \regep/data_out_buffer_reg[27]  ( .D(alutwo_out[27]), .E(n1986), 
        .CK(clk), .Q(regep_out[27]) );
  EDFFX1TS \regep/data_out_buffer_reg[28]  ( .D(alutwo_out[28]), .E(n1986), 
        .CK(clk), .Q(regep_out[28]) );
  EDFFX1TS \regep/data_out_buffer_reg[29]  ( .D(alutwo_out[29]), .E(n1986), 
        .CK(clk), .Q(regep_out[29]) );
  EDFFX1TS \regep/data_out_buffer_reg[30]  ( .D(alutwo_out[30]), .E(n1986), 
        .CK(clk), .Q(regep_out[30]) );
  EDFFX1TS \regep/data_out_buffer_reg[31]  ( .D(alutwo_out[31]), .E(n1986), 
        .CK(clk), .Q(regep_out[31]) );
  EDFFX1TS \regeq/data_out_buffer_reg[0]  ( .D(alutwo_out[0]), .E(n1988), .CK(
        clk), .Q(regeq_out[0]) );
  EDFFX1TS \regeq/data_out_buffer_reg[1]  ( .D(alutwo_out[1]), .E(n1988), .CK(
        clk), .Q(regeq_out[1]) );
  EDFFX1TS \regeq/data_out_buffer_reg[2]  ( .D(alutwo_out[2]), .E(n1988), .CK(
        clk), .Q(regeq_out[2]) );
  EDFFX1TS \regeq/data_out_buffer_reg[3]  ( .D(alutwo_out[3]), .E(n1988), .CK(
        clk), .Q(regeq_out[3]) );
  EDFFX1TS \regeq/data_out_buffer_reg[4]  ( .D(alutwo_out[4]), .E(n1988), .CK(
        clk), .Q(regeq_out[4]) );
  EDFFX1TS \regeq/data_out_buffer_reg[5]  ( .D(alutwo_out[5]), .E(n1988), .CK(
        clk), .Q(regeq_out[5]) );
  EDFFX1TS \regeq/data_out_buffer_reg[6]  ( .D(alutwo_out[6]), .E(n1988), .CK(
        clk), .Q(regeq_out[6]) );
  EDFFX1TS \regeq/data_out_buffer_reg[7]  ( .D(alutwo_out[7]), .E(n1988), .CK(
        clk), .Q(regeq_out[7]) );
  EDFFX1TS \regeq/data_out_buffer_reg[8]  ( .D(alutwo_out[8]), .E(n1988), .CK(
        clk), .Q(regeq_out[8]) );
  EDFFX1TS \regeq/data_out_buffer_reg[9]  ( .D(alutwo_out[9]), .E(n1988), .CK(
        clk), .Q(regeq_out[9]) );
  EDFFX1TS \regeq/data_out_buffer_reg[10]  ( .D(alutwo_out[10]), .E(n1988), 
        .CK(clk), .Q(regeq_out[10]) );
  EDFFX1TS \regeq/data_out_buffer_reg[11]  ( .D(alutwo_out[11]), .E(n1988), 
        .CK(clk), .Q(regeq_out[11]) );
  EDFFX1TS \regeq/data_out_buffer_reg[12]  ( .D(alutwo_out[12]), .E(n1988), 
        .CK(clk), .Q(regeq_out[12]) );
  EDFFX1TS \regeq/data_out_buffer_reg[13]  ( .D(alutwo_out[13]), .E(n1988), 
        .CK(clk), .Q(regeq_out[13]) );
  EDFFX1TS \regeq/data_out_buffer_reg[14]  ( .D(alutwo_out[14]), .E(n1988), 
        .CK(clk), .Q(regeq_out[14]) );
  EDFFX1TS \regeq/data_out_buffer_reg[15]  ( .D(alutwo_out[15]), .E(n1988), 
        .CK(clk), .Q(regeq_out[15]) );
  EDFFX1TS \regeq/data_out_buffer_reg[16]  ( .D(alutwo_out[16]), .E(n1988), 
        .CK(clk), .Q(regeq_out[16]) );
  EDFFX1TS \regeq/data_out_buffer_reg[17]  ( .D(alutwo_out[17]), .E(n1988), 
        .CK(clk), .Q(regeq_out[17]) );
  EDFFX1TS \regeq/data_out_buffer_reg[18]  ( .D(alutwo_out[18]), .E(n1988), 
        .CK(clk), .Q(regeq_out[18]) );
  EDFFX1TS \regeq/data_out_buffer_reg[19]  ( .D(alutwo_out[19]), .E(n1988), 
        .CK(clk), .Q(regeq_out[19]) );
  EDFFX1TS \regeq/data_out_buffer_reg[20]  ( .D(alutwo_out[20]), .E(n1988), 
        .CK(clk), .Q(regeq_out[20]) );
  EDFFX1TS \regeq/data_out_buffer_reg[21]  ( .D(alutwo_out[21]), .E(n1988), 
        .CK(clk), .Q(regeq_out[21]) );
  EDFFX1TS \regeq/data_out_buffer_reg[22]  ( .D(alutwo_out[22]), .E(n1988), 
        .CK(clk), .Q(regeq_out[22]) );
  EDFFX1TS \regeq/data_out_buffer_reg[23]  ( .D(alutwo_out[23]), .E(n1988), 
        .CK(clk), .Q(regeq_out[23]) );
  EDFFX1TS \regeq/data_out_buffer_reg[24]  ( .D(alutwo_out[24]), .E(n1988), 
        .CK(clk), .Q(regeq_out[24]) );
  EDFFX1TS \regeq/data_out_buffer_reg[25]  ( .D(alutwo_out[25]), .E(n1988), 
        .CK(clk), .Q(regeq_out[25]) );
  EDFFX1TS \regeq/data_out_buffer_reg[26]  ( .D(alutwo_out[26]), .E(n1988), 
        .CK(clk), .Q(regeq_out[26]) );
  EDFFX1TS \regeq/data_out_buffer_reg[27]  ( .D(alutwo_out[27]), .E(n1988), 
        .CK(clk), .Q(regeq_out[27]) );
  EDFFX1TS \regeq/data_out_buffer_reg[28]  ( .D(alutwo_out[28]), .E(n1988), 
        .CK(clk), .Q(regeq_out[28]) );
  EDFFX1TS \regeq/data_out_buffer_reg[29]  ( .D(alutwo_out[29]), .E(n1988), 
        .CK(clk), .Q(regeq_out[29]) );
  EDFFX1TS \regeq/data_out_buffer_reg[30]  ( .D(alutwo_out[30]), .E(n1988), 
        .CK(clk), .Q(regeq_out[30]) );
  EDFFX1TS \regeq/data_out_buffer_reg[31]  ( .D(alutwo_out[31]), .E(n1988), 
        .CK(clk), .Q(regeq_out[31]) );
  EDFFX1TS \regr/data_out_buffer_reg[0]  ( .D(aluone_out[0]), .E(n1993), .CK(
        clk), .Q(regr_out[0]) );
  EDFFX1TS \regr/data_out_buffer_reg[1]  ( .D(aluone_out[1]), .E(n1993), .CK(
        clk), .Q(regr_out[1]) );
  EDFFX1TS \regr/data_out_buffer_reg[2]  ( .D(aluone_out[2]), .E(n1993), .CK(
        clk), .Q(regr_out[2]) );
  EDFFX1TS \regr/data_out_buffer_reg[3]  ( .D(aluone_out[3]), .E(n1993), .CK(
        clk), .Q(regr_out[3]) );
  EDFFX1TS \regr/data_out_buffer_reg[4]  ( .D(aluone_out[4]), .E(n1993), .CK(
        clk), .Q(regr_out[4]) );
  EDFFX1TS \regr/data_out_buffer_reg[5]  ( .D(aluone_out[5]), .E(n1993), .CK(
        clk), .Q(regr_out[5]) );
  EDFFX1TS \regr/data_out_buffer_reg[6]  ( .D(aluone_out[6]), .E(n1993), .CK(
        clk), .Q(regr_out[6]) );
  EDFFX1TS \regr/data_out_buffer_reg[7]  ( .D(aluone_out[7]), .E(n1993), .CK(
        clk), .Q(regr_out[7]) );
  EDFFX1TS \regr/data_out_buffer_reg[8]  ( .D(aluone_out[8]), .E(n1993), .CK(
        clk), .Q(regr_out[8]) );
  EDFFX1TS \regr/data_out_buffer_reg[9]  ( .D(aluone_out[9]), .E(n1993), .CK(
        clk), .Q(regr_out[9]) );
  EDFFX1TS \regr/data_out_buffer_reg[10]  ( .D(aluone_out[10]), .E(n1993), 
        .CK(clk), .Q(regr_out[10]) );
  EDFFX1TS \regr/data_out_buffer_reg[11]  ( .D(aluone_out[11]), .E(n1993), 
        .CK(clk), .Q(regr_out[11]) );
  EDFFX1TS \regr/data_out_buffer_reg[12]  ( .D(aluone_out[12]), .E(n1993), 
        .CK(clk), .Q(regr_out[12]) );
  EDFFX1TS \regr/data_out_buffer_reg[13]  ( .D(aluone_out[13]), .E(n1993), 
        .CK(clk), .Q(regr_out[13]) );
  EDFFX1TS \regr/data_out_buffer_reg[14]  ( .D(aluone_out[14]), .E(n1993), 
        .CK(clk), .Q(regr_out[14]) );
  EDFFX1TS \regr/data_out_buffer_reg[15]  ( .D(aluone_out[15]), .E(n1993), 
        .CK(clk), .Q(regr_out[15]) );
  EDFFX1TS \regr/data_out_buffer_reg[16]  ( .D(aluone_out[16]), .E(n1993), 
        .CK(clk), .Q(regr_out[16]) );
  EDFFX1TS \regr/data_out_buffer_reg[17]  ( .D(aluone_out[17]), .E(n1993), 
        .CK(clk), .Q(regr_out[17]) );
  EDFFX1TS \regr/data_out_buffer_reg[18]  ( .D(aluone_out[18]), .E(n1993), 
        .CK(clk), .Q(regr_out[18]) );
  EDFFX1TS \regr/data_out_buffer_reg[19]  ( .D(aluone_out[19]), .E(n1993), 
        .CK(clk), .Q(regr_out[19]) );
  EDFFX1TS \regr/data_out_buffer_reg[20]  ( .D(aluone_out[20]), .E(n1993), 
        .CK(clk), .Q(regr_out[20]) );
  EDFFX1TS \regr/data_out_buffer_reg[21]  ( .D(aluone_out[21]), .E(n1993), 
        .CK(clk), .Q(regr_out[21]) );
  EDFFX1TS \regr/data_out_buffer_reg[22]  ( .D(aluone_out[22]), .E(n1993), 
        .CK(clk), .Q(regr_out[22]) );
  EDFFX1TS \regr/data_out_buffer_reg[23]  ( .D(aluone_out[23]), .E(n1993), 
        .CK(clk), .Q(regr_out[23]) );
  EDFFX1TS \regr/data_out_buffer_reg[24]  ( .D(aluone_out[24]), .E(n1993), 
        .CK(clk), .Q(regr_out[24]) );
  EDFFX1TS \regr/data_out_buffer_reg[25]  ( .D(aluone_out[25]), .E(n1993), 
        .CK(clk), .Q(regr_out[25]) );
  EDFFX1TS \regr/data_out_buffer_reg[26]  ( .D(aluone_out[26]), .E(n1993), 
        .CK(clk), .Q(regr_out[26]) );
  EDFFX1TS \regr/data_out_buffer_reg[27]  ( .D(aluone_out[27]), .E(n1993), 
        .CK(clk), .Q(regr_out[27]) );
  EDFFX1TS \regr/data_out_buffer_reg[28]  ( .D(aluone_out[28]), .E(n1993), 
        .CK(clk), .Q(regr_out[28]) );
  EDFFX1TS \regr/data_out_buffer_reg[29]  ( .D(aluone_out[29]), .E(n1993), 
        .CK(clk), .Q(regr_out[29]) );
  EDFFX1TS \regr/data_out_buffer_reg[30]  ( .D(aluone_out[30]), .E(n1993), 
        .CK(clk), .Q(regr_out[30]) );
  EDFFX1TS \regr/data_out_buffer_reg[31]  ( .D(aluone_out[31]), .E(n1993), 
        .CK(clk), .Q(regr_out[31]) );
  EDFFX1TS \regindex/data_out_buffer_reg[0]  ( .D(m13_out[0]), .E(reg_index), 
        .CK(clk), .Q(regindex_out[0]) );
  EDFFX1TS \regindex/data_out_buffer_reg[1]  ( .D(m13_out[1]), .E(reg_index), 
        .CK(clk), .Q(regindex_out[1]) );
  EDFFX1TS \regindex/data_out_buffer_reg[2]  ( .D(m13_out[2]), .E(reg_index), 
        .CK(clk), .Q(regindex_out[2]) );
  EDFFX1TS \regindex/data_out_buffer_reg[3]  ( .D(m13_out[3]), .E(reg_index), 
        .CK(clk), .QN(n4773) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[0]  ( .D(m3_out[0]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[0]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[1]  ( .D(m3_out[1]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[1]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[2]  ( .D(m3_out[2]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[2]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[3]  ( .D(m3_out[3]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[3]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[4]  ( .D(m3_out[4]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[4]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[5]  ( .D(m3_out[5]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[5]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[6]  ( .D(m3_out[6]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[6]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[7]  ( .D(m3_out[7]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[7]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[8]  ( .D(m3_out[8]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[8]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[9]  ( .D(m3_out[9]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[9]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[10]  ( .D(m3_out[10]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[10]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[11]  ( .D(m3_out[11]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[11]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[12]  ( .D(m3_out[12]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[12]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[13]  ( .D(m3_out[13]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[13]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[14]  ( .D(m3_out[14]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[14]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[15]  ( .D(m3_out[15]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[15]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[16]  ( .D(m3_out[16]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[16]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[17]  ( .D(m3_out[17]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[17]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[18]  ( .D(m3_out[18]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[18]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[19]  ( .D(m3_out[19]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[19]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[21]  ( .D(m3_out[21]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[21]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[22]  ( .D(m3_out[22]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[22]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[23]  ( .D(m3_out[23]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[23]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[24]  ( .D(m3_out[24]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[24]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[28]  ( .D(m3_out[28]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[28]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[30]  ( .D(m3_out[30]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[30]) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[31]  ( .D(m3_out[31]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[31]) );
  EDFFX1TS \regsum/data_out_buffer_reg[4]  ( .D(m2_out[4]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[4]) );
  EDFFX1TS \regsum/data_out_buffer_reg[8]  ( .D(m2_out[8]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[8]) );
  EDFFX1TS \regsum/data_out_buffer_reg[9]  ( .D(m2_out[9]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[9]) );
  EDFFX1TS \regsum/data_out_buffer_reg[14]  ( .D(m2_out[14]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[14]) );
  EDFFX1TS \regsum/data_out_buffer_reg[16]  ( .D(m2_out[16]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[16]) );
  EDFFX1TS \regsum/data_out_buffer_reg[19]  ( .D(m2_out[19]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[19]) );
  EDFFX1TS \regsum/data_out_buffer_reg[27]  ( .D(m2_out[27]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[27]) );
  EDFFX1TS \regsum/data_out_buffer_reg[31]  ( .D(m2_out[31]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[31]) );
  EDFFX1TS \regmb/data_out_buffer_reg[0]  ( .D(rf_bout[0]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[0]) );
  EDFFX1TS \regmb/data_out_buffer_reg[1]  ( .D(rf_bout[1]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[1]) );
  EDFFX1TS \regmb/data_out_buffer_reg[2]  ( .D(rf_bout[2]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[2]) );
  EDFFX1TS \regmb/data_out_buffer_reg[3]  ( .D(rf_bout[3]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[3]) );
  EDFFX1TS \regmb/data_out_buffer_reg[4]  ( .D(rf_bout[4]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[4]) );
  EDFFX1TS \regmb/data_out_buffer_reg[5]  ( .D(rf_bout[5]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[5]) );
  EDFFX1TS \regmb/data_out_buffer_reg[6]  ( .D(rf_bout[6]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[6]) );
  EDFFX1TS \regmb/data_out_buffer_reg[7]  ( .D(rf_bout[7]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[7]) );
  EDFFX1TS \regmb/data_out_buffer_reg[8]  ( .D(rf_bout[8]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[8]) );
  EDFFX1TS \regmb/data_out_buffer_reg[9]  ( .D(rf_bout[9]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[9]) );
  EDFFX1TS \regeb/data_out_buffer_reg[0]  ( .D(rf_bout[23]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[0]) );
  EDFFX1TS \regeb/data_out_buffer_reg[1]  ( .D(rf_bout[24]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[1]) );
  EDFFX1TS \regeb/data_out_buffer_reg[2]  ( .D(rf_bout[25]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[2]) );
  EDFFX1TS \regeb/data_out_buffer_reg[3]  ( .D(rf_bout[26]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[3]) );
  EDFFX1TS \regeb/data_out_buffer_reg[4]  ( .D(rf_bout[27]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[4]) );
  EDFFX1TS \regeb/data_out_buffer_reg[5]  ( .D(rf_bout[28]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[5]) );
  EDFFX1TS \regeb/data_out_buffer_reg[6]  ( .D(rf_bout[29]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[6]) );
  EDFFX1TS \regeb/data_out_buffer_reg[7]  ( .D(rf_bout[30]), .E(reg_eb), .CK(
        clk), .Q(regeb_out[7]) );
  EDFFX1TS \regsb/data_out_buffer_reg  ( .D(rf_bout[31]), .E(reg_sb), .CK(clk), 
        .Q(regsb_out) );
  EDFFX1TS \regmc/data_out_buffer_reg[0]  ( .D(rf_aout[0]), .E(n1990), .CK(clk), .Q(regmc_out[0]) );
  EDFFX1TS \regmc/data_out_buffer_reg[1]  ( .D(rf_aout[1]), .E(n1990), .CK(clk), .Q(regmc_out[1]) );
  EDFFX1TS \regmc/data_out_buffer_reg[2]  ( .D(rf_aout[2]), .E(n1990), .CK(clk), .Q(regmc_out[2]) );
  EDFFX1TS \regmc/data_out_buffer_reg[3]  ( .D(rf_aout[3]), .E(n1990), .CK(clk), .Q(regmc_out[3]) );
  EDFFX1TS \regmc/data_out_buffer_reg[4]  ( .D(rf_aout[4]), .E(n1990), .CK(clk), .Q(regmc_out[4]) );
  EDFFX1TS \regmc/data_out_buffer_reg[5]  ( .D(rf_aout[5]), .E(n1990), .CK(clk), .Q(regmc_out[5]) );
  EDFFX1TS \regmc/data_out_buffer_reg[6]  ( .D(rf_aout[6]), .E(n1990), .CK(clk), .Q(regmc_out[6]) );
  EDFFX1TS \regmc/data_out_buffer_reg[7]  ( .D(rf_aout[7]), .E(n1990), .CK(clk), .Q(regmc_out[7]) );
  EDFFX1TS \regmc/data_out_buffer_reg[8]  ( .D(rf_aout[8]), .E(n1990), .CK(clk), .Q(regmc_out[8]) );
  EDFFX1TS \regmc/data_out_buffer_reg[9]  ( .D(rf_aout[9]), .E(n1990), .CK(clk), .Q(regmc_out[9]) );
  EDFFX1TS \regmc/data_out_buffer_reg[10]  ( .D(rf_aout[10]), .E(n1990), .CK(
        clk), .Q(regmc_out[10]) );
  EDFFX1TS \regmc/data_out_buffer_reg[11]  ( .D(rf_aout[11]), .E(n1990), .CK(
        clk), .Q(regmc_out[11]) );
  EDFFX1TS \regmc/data_out_buffer_reg[12]  ( .D(rf_aout[12]), .E(n1990), .CK(
        clk), .Q(regmc_out[12]) );
  EDFFX1TS \regmc/data_out_buffer_reg[13]  ( .D(rf_aout[13]), .E(n1990), .CK(
        clk), .Q(regmc_out[13]) );
  EDFFX1TS \regmc/data_out_buffer_reg[14]  ( .D(rf_aout[14]), .E(n1990), .CK(
        clk), .Q(regmc_out[14]) );
  EDFFX1TS \regmc/data_out_buffer_reg[15]  ( .D(rf_aout[15]), .E(n1990), .CK(
        clk), .Q(regmc_out[15]) );
  EDFFX1TS \regmc/data_out_buffer_reg[16]  ( .D(rf_aout[16]), .E(n1990), .CK(
        clk), .Q(regmc_out[16]) );
  EDFFX1TS \regmc/data_out_buffer_reg[17]  ( .D(rf_aout[17]), .E(n1990), .CK(
        clk), .Q(regmc_out[17]) );
  EDFFX1TS \regmc/data_out_buffer_reg[18]  ( .D(rf_aout[18]), .E(n1990), .CK(
        clk), .Q(regmc_out[18]) );
  EDFFX1TS \regmc/data_out_buffer_reg[19]  ( .D(rf_aout[19]), .E(n1990), .CK(
        clk), .Q(regmc_out[19]) );
  EDFFX1TS \regmc/data_out_buffer_reg[20]  ( .D(rf_aout[20]), .E(n1990), .CK(
        clk), .Q(regmc_out[20]) );
  EDFFX1TS \regmc/data_out_buffer_reg[21]  ( .D(rf_aout[21]), .E(n1990), .CK(
        clk), .Q(regmc_out[21]) );
  EDFFX1TS \regmc/data_out_buffer_reg[22]  ( .D(rf_aout[22]), .E(n1990), .CK(
        clk), .Q(regmc_out[22]) );
  EDFFX1TS \regec/data_out_buffer_reg[0]  ( .D(rf_aout[23]), .E(reg_ec), .CK(
        clk), .Q(regec_out[0]) );
  EDFFX1TS \regec/data_out_buffer_reg[1]  ( .D(rf_aout[24]), .E(reg_ec), .CK(
        clk), .Q(regec_out[1]) );
  EDFFX1TS \regec/data_out_buffer_reg[2]  ( .D(rf_aout[25]), .E(reg_ec), .CK(
        clk), .Q(regec_out[2]) );
  EDFFX1TS \regec/data_out_buffer_reg[3]  ( .D(rf_aout[26]), .E(reg_ec), .CK(
        clk), .Q(regec_out[3]) );
  EDFFX1TS \regec/data_out_buffer_reg[4]  ( .D(rf_aout[27]), .E(reg_ec), .CK(
        clk), .Q(regec_out[4]) );
  EDFFX1TS \regec/data_out_buffer_reg[5]  ( .D(rf_aout[28]), .E(reg_ec), .CK(
        clk), .Q(regec_out[5]) );
  EDFFX1TS \regec/data_out_buffer_reg[6]  ( .D(rf_aout[29]), .E(reg_ec), .CK(
        clk), .Q(regec_out[6]) );
  EDFFX1TS \regec/data_out_buffer_reg[7]  ( .D(rf_aout[30]), .E(reg_ec), .CK(
        clk), .Q(regec_out[7]) );
  EDFFX1TS \regsc/data_out_buffer_reg  ( .D(rf_aout[31]), .E(reg_sc), .CK(clk), 
        .Q(regsc_out) );
  EDFFX1TS \regms/data_out_buffer_reg[0]  ( .D(m4_out[0]), .E(n1989), .CK(clk), 
        .Q(regms_out[0]) );
  EDFFX1TS \regms/data_out_buffer_reg[1]  ( .D(m4_out[1]), .E(n1989), .CK(clk), 
        .Q(regms_out[1]) );
  EDFFX1TS \regms/data_out_buffer_reg[2]  ( .D(m4_out[2]), .E(n1989), .CK(clk), 
        .Q(regms_out[2]) );
  EDFFX1TS \regms/data_out_buffer_reg[3]  ( .D(m4_out[3]), .E(n1989), .CK(clk), 
        .Q(regms_out[3]) );
  EDFFX1TS \regms/data_out_buffer_reg[4]  ( .D(m4_out[4]), .E(n1989), .CK(clk), 
        .Q(regms_out[4]) );
  EDFFX1TS \regms/data_out_buffer_reg[5]  ( .D(m4_out[5]), .E(n1989), .CK(clk), 
        .Q(regms_out[5]) );
  EDFFX1TS \regms/data_out_buffer_reg[6]  ( .D(m4_out[6]), .E(n1989), .CK(clk), 
        .Q(regms_out[6]) );
  EDFFX1TS \regms/data_out_buffer_reg[7]  ( .D(m4_out[7]), .E(n1989), .CK(clk), 
        .Q(regms_out[7]) );
  EDFFX1TS \regms/data_out_buffer_reg[8]  ( .D(m4_out[8]), .E(n1989), .CK(clk), 
        .Q(regms_out[8]) );
  EDFFX1TS \regms/data_out_buffer_reg[9]  ( .D(m4_out[9]), .E(n1989), .CK(clk), 
        .Q(regms_out[9]) );
  EDFFX1TS \regms/data_out_buffer_reg[10]  ( .D(m4_out[10]), .E(n1989), .CK(
        clk), .Q(regms_out[10]) );
  EDFFX1TS \regms/data_out_buffer_reg[11]  ( .D(m4_out[11]), .E(n1989), .CK(
        clk), .Q(regms_out[11]) );
  EDFFX1TS \regms/data_out_buffer_reg[12]  ( .D(m4_out[12]), .E(n1989), .CK(
        clk), .Q(regms_out[12]) );
  EDFFX1TS \regms/data_out_buffer_reg[13]  ( .D(m4_out[13]), .E(n1989), .CK(
        clk), .Q(regms_out[13]) );
  EDFFX1TS \regms/data_out_buffer_reg[14]  ( .D(m4_out[14]), .E(n1989), .CK(
        clk), .Q(regms_out[14]) );
  EDFFX1TS \regms/data_out_buffer_reg[15]  ( .D(m4_out[15]), .E(n1989), .CK(
        clk), .Q(regms_out[15]) );
  EDFFX1TS \regms/data_out_buffer_reg[16]  ( .D(m4_out[16]), .E(n1989), .CK(
        clk), .Q(regms_out[16]) );
  EDFFX1TS \regms/data_out_buffer_reg[17]  ( .D(m4_out[17]), .E(n1989), .CK(
        clk), .Q(regms_out[17]) );
  EDFFX1TS \regms/data_out_buffer_reg[18]  ( .D(m4_out[18]), .E(n1989), .CK(
        clk), .Q(regms_out[18]) );
  EDFFX1TS \regms/data_out_buffer_reg[19]  ( .D(m4_out[19]), .E(n1989), .CK(
        clk), .Q(regms_out[19]) );
  EDFFX1TS \regms/data_out_buffer_reg[20]  ( .D(m4_out[20]), .E(n1989), .CK(
        clk), .Q(regms_out[20]) );
  EDFFX1TS \regms/data_out_buffer_reg[21]  ( .D(m4_out[21]), .E(n1989), .CK(
        clk), .Q(regms_out[21]) );
  EDFFX1TS \regms/data_out_buffer_reg[22]  ( .D(m4_out[22]), .E(n1989), .CK(
        clk), .Q(regms_out[22]) );
  EDFFX1TS \regms/data_out_buffer_reg[23]  ( .D(m4_out[23]), .E(n1989), .CK(
        clk), .Q(regms_out[23]) );
  EDFFX1TS \regms/data_out_buffer_reg[24]  ( .D(m4_out[24]), .E(n1989), .CK(
        clk), .Q(regms_out[24]) );
  EDFFX1TS \regms/data_out_buffer_reg[25]  ( .D(m4_out[25]), .E(n1989), .CK(
        clk), .Q(regms_out[25]) );
  EDFFX1TS \regms/data_out_buffer_reg[26]  ( .D(m4_out[26]), .E(n1989), .CK(
        clk), .Q(regms_out[26]) );
  EDFFX1TS \regms/data_out_buffer_reg[27]  ( .D(m4_out[27]), .E(n1989), .CK(
        clk), .Q(regms_out[27]) );
  EDFFX1TS \regms/data_out_buffer_reg[28]  ( .D(m4_out[28]), .E(n1989), .CK(
        clk), .Q(regms_out[28]) );
  EDFFX1TS \regms/data_out_buffer_reg[29]  ( .D(m4_out[29]), .E(n1989), .CK(
        clk), .Q(n4821) );
  EDFFX1TS \regms/data_out_buffer_reg[30]  ( .D(m4_out[30]), .E(n1989), .CK(
        clk), .Q(regms_out[30]) );
  EDFFX1TS \regms/data_out_buffer_reg[31]  ( .D(m4_out[31]), .E(n1989), .CK(
        clk), .Q(regms_out[31]) );
  DFFQX1TS \ssrms0/tmp_reg[9]  ( .D(n1888), .CK(clk), .Q(ssrms0_out[9]) );
  TLATXLTS \alutwo/Cout_reg  ( .G(\alutwo/N324 ), .D(\alutwo/N325 ), .Q(
        Couttwo) );
  TLATXLTS \aluone/Cout_reg  ( .G(\aluone/N324 ), .D(\aluone/N325 ), .Q(
        Coutone) );
  DFFQX1TS \srmp/tmp_reg[61]  ( .D(n1876), .CK(clk), .Q(srmp_out[61]) );
  DFFQX1TS \srmp/tmp_reg[59]  ( .D(n1874), .CK(clk), .Q(srmp_out[59]) );
  DFFQX1TS \srmp/tmp_reg[57]  ( .D(n1872), .CK(clk), .Q(srmp_out[57]) );
  DFFQX1TS \srmp/tmp_reg[55]  ( .D(n1870), .CK(clk), .Q(srmp_out[55]) );
  DFFQX1TS \srmp/tmp_reg[63]  ( .D(n1878), .CK(clk), .Q(srmp_out[63]) );
  DFFQX1TS \srmp/tmp_reg[53]  ( .D(n1868), .CK(clk), .Q(srmp_out[53]) );
  DFFQX1TS \srmp/tmp_reg[49]  ( .D(n1864), .CK(clk), .Q(srmp_out[49]) );
  DFFQX1TS \srmp/tmp_reg[46]  ( .D(n1861), .CK(clk), .Q(srmp_out[46]) );
  DFFQX1TS \srmp/tmp_reg[9]  ( .D(n1824), .CK(clk), .Q(srmp_out[9]) );
  DFFQX1TS \srmp/tmp_reg[4]  ( .D(n1819), .CK(clk), .Q(srmp_out[4]) );
  DFFQX1TS \srmp/tmp_reg[51]  ( .D(n1866), .CK(clk), .Q(srmp_out[51]) );
  DFFQX1TS \srmp/tmp_reg[50]  ( .D(n1865), .CK(clk), .Q(srmp_out[50]) );
  DFFQX1TS \srmp/tmp_reg[22]  ( .D(n1837), .CK(clk), .Q(srmp_out[22]) );
  DFFQX1TS \srmp/tmp_reg[21]  ( .D(n1836), .CK(clk), .Q(srmp_out[21]) );
  DFFQX1TS \srmp/tmp_reg[20]  ( .D(n1835), .CK(clk), .Q(srmp_out[20]) );
  DFFQX1TS \srmp/tmp_reg[19]  ( .D(n1834), .CK(clk), .Q(srmp_out[19]) );
  DFFQX1TS \srmp/tmp_reg[17]  ( .D(n1832), .CK(clk), .Q(srmp_out[17]) );
  DFFQX1TS \srmp/tmp_reg[16]  ( .D(n1831), .CK(clk), .Q(srmp_out[16]) );
  DFFQX1TS \srmp/tmp_reg[15]  ( .D(n1830), .CK(clk), .Q(srmp_out[15]) );
  DFFQX1TS \srmp/tmp_reg[14]  ( .D(n1829), .CK(clk), .Q(srmp_out[14]) );
  DFFQX1TS \srmp/tmp_reg[13]  ( .D(n1828), .CK(clk), .Q(srmp_out[13]) );
  DFFQX1TS \srmp/tmp_reg[12]  ( .D(n1827), .CK(clk), .Q(srmp_out[12]) );
  DFFQX1TS \srmp/tmp_reg[11]  ( .D(n1826), .CK(clk), .Q(srmp_out[11]) );
  DFFQX1TS \srmp/tmp_reg[10]  ( .D(n1825), .CK(clk), .Q(srmp_out[10]) );
  DFFQX1TS \srmp/tmp_reg[7]  ( .D(n1822), .CK(clk), .Q(srmp_out[7]) );
  DFFQX1TS \srmp/tmp_reg[6]  ( .D(n1821), .CK(clk), .Q(srmp_out[6]) );
  DFFQX1TS \srmp/tmp_reg[5]  ( .D(n1820), .CK(clk), .Q(srmp_out[5]) );
  DFFQX1TS \srmp/tmp_reg[3]  ( .D(n1818), .CK(clk), .Q(srmp_out[3]) );
  DFFQX1TS \srmp/tmp_reg[62]  ( .D(n1877), .CK(clk), .Q(srmp_out[62]) );
  DFFQX1TS \srmp/tmp_reg[60]  ( .D(n1875), .CK(clk), .Q(srmp_out[60]) );
  DFFQX1TS \srmp/tmp_reg[58]  ( .D(n1873), .CK(clk), .Q(srmp_out[58]) );
  DFFQX1TS \srmp/tmp_reg[56]  ( .D(n1871), .CK(clk), .Q(srmp_out[56]) );
  DFFQX1TS \srmp/tmp_reg[54]  ( .D(n1869), .CK(clk), .Q(srmp_out[54]) );
  DFFQX1TS \srmp/tmp_reg[52]  ( .D(n1867), .CK(clk), .Q(srmp_out[52]) );
  DFFQX1TS \srmp/tmp_reg[48]  ( .D(n1863), .CK(clk), .Q(srmp_out[48]) );
  DFFQX1TS \srmp/tmp_reg[18]  ( .D(n1833), .CK(clk), .Q(srmp_out[18]) );
  DFFQX1TS \srmp/tmp_reg[8]  ( .D(n1823), .CK(clk), .Q(srmp_out[8]) );
  DFFQX1TS \srmp/tmp_reg[2]  ( .D(n1817), .CK(clk), .Q(srmp_out[2]) );
  DFFQX1TS \srmp/tmp_reg[47]  ( .D(n1862), .CK(clk), .Q(srmp_out[47]) );
  DFFQX1TS \regsp/data_out_buffer_reg  ( .D(n1683), .CK(clk), .Q(regsp_out) );
  DFFQX1TS \srmp/tmp_reg[0]  ( .D(n1815), .CK(clk), .Q(srmp_out[0]) );
  DFFQX1TS \srmp/tmp_reg[1]  ( .D(n1816), .CK(clk), .Q(srmp_out[1]) );
  DFFQX1TS \srmp/tmp_reg[44]  ( .D(n1859), .CK(clk), .Q(srmp_out[44]) );
  DFFQX1TS \srmp/tmp_reg[39]  ( .D(n1854), .CK(clk), .Q(srmp_out[39]) );
  DFFQX1TS \srmp/tmp_reg[33]  ( .D(n1848), .CK(clk), .Q(srmp_out[33]) );
  DFFQX1TS \srmp/tmp_reg[31]  ( .D(n1846), .CK(clk), .Q(srmp_out[31]) );
  DFFQX1TS \srmp/tmp_reg[27]  ( .D(n1842), .CK(clk), .Q(srmp_out[27]) );
  DFFQX1TS \srmp/tmp_reg[24]  ( .D(n1839), .CK(clk), .Q(srmp_out[24]) );
  DFFQX1TS \srmp/tmp_reg[43]  ( .D(n1858), .CK(clk), .Q(srmp_out[43]) );
  DFFQX1TS \srmp/tmp_reg[41]  ( .D(n1856), .CK(clk), .Q(srmp_out[41]) );
  DFFQX1TS \srmp/tmp_reg[40]  ( .D(n1855), .CK(clk), .Q(srmp_out[40]) );
  DFFQX1TS \srmp/tmp_reg[38]  ( .D(n1853), .CK(clk), .Q(srmp_out[38]) );
  DFFQX1TS \srmp/tmp_reg[36]  ( .D(n1851), .CK(clk), .Q(srmp_out[36]) );
  DFFQX1TS \srmp/tmp_reg[35]  ( .D(n1850), .CK(clk), .Q(srmp_out[35]) );
  DFFQX1TS \srmp/tmp_reg[34]  ( .D(n1849), .CK(clk), .Q(srmp_out[34]) );
  DFFQX1TS \srmp/tmp_reg[29]  ( .D(n1844), .CK(clk), .Q(srmp_out[29]) );
  DFFQX1TS \srmp/tmp_reg[28]  ( .D(n1843), .CK(clk), .Q(srmp_out[28]) );
  DFFQX1TS \srmp/tmp_reg[25]  ( .D(n1840), .CK(clk), .Q(srmp_out[25]) );
  DFFQX1TS \srmp/tmp_reg[23]  ( .D(n1838), .CK(clk), .Q(srmp_out[23]) );
  DFFQX1TS \srmp/tmp_reg[45]  ( .D(n1860), .CK(clk), .Q(srmp_out[45]) );
  DFFQX1TS \srmp/tmp_reg[42]  ( .D(n1857), .CK(clk), .Q(srmp_out[42]) );
  DFFQX1TS \srmp/tmp_reg[37]  ( .D(n1852), .CK(clk), .Q(srmp_out[37]) );
  DFFQX1TS \srmp/tmp_reg[32]  ( .D(n1847), .CK(clk), .Q(srmp_out[32]) );
  DFFQX1TS \srmp/tmp_reg[30]  ( .D(n1845), .CK(clk), .Q(srmp_out[30]) );
  DFFQX1TS \srmp/tmp_reg[26]  ( .D(n1841), .CK(clk), .Q(srmp_out[26]) );
  DFFQX1TS \count/data_out_reg[4]  ( .D(n4779), .CK(clk), .Q(count_out[4]) );
  DFFQX1TS \count/data_out_reg[5]  ( .D(\count/N34 ), .CK(clk), .Q(
        count_out[5]) );
  DFFQX1TS \count/data_out_reg[2]  ( .D(n4780), .CK(clk), .Q(count_out[2]) );
  DFFQX1TS \count/data_out_reg[3]  ( .D(\count/N32 ), .CK(clk), .Q(
        count_out[3]) );
  DFFQX1TS \srmq/tmp_reg[61]  ( .D(n1780), .CK(clk), .Q(srmq_out[61]) );
  DFFQX1TS \regsq/data_out_buffer_reg  ( .D(n1682), .CK(clk), .Q(regsq_out) );
  DFFQX1TS \ssrms0/tmp_reg[40]  ( .D(n1919), .CK(clk), .Q(ssrms0_out[40]) );
  DFFQX1TS \ssrms0/tmp_reg[61]  ( .D(n1940), .CK(clk), .Q(ssrms0_out[61]) );
  DFFQX1TS \ssrms0/tmp_reg[59]  ( .D(n1938), .CK(clk), .Q(ssrms0_out[59]) );
  DFFQX1TS \ssrms0/tmp_reg[57]  ( .D(n1936), .CK(clk), .Q(ssrms0_out[57]) );
  DFFQX1TS \ssrms0/tmp_reg[55]  ( .D(n1934), .CK(clk), .Q(ssrms0_out[55]) );
  DFFQX1TS \ssrms0/tmp_reg[53]  ( .D(n1932), .CK(clk), .Q(ssrms0_out[53]) );
  DFFQX1TS \ssrms0/tmp_reg[51]  ( .D(n1930), .CK(clk), .Q(ssrms0_out[51]) );
  DFFQX1TS \ssrms0/tmp_reg[49]  ( .D(n1928), .CK(clk), .Q(ssrms0_out[49]) );
  DFFQX1TS \ssrms0/tmp_reg[47]  ( .D(n1926), .CK(clk), .Q(ssrms0_out[47]) );
  DFFQX1TS \ssrms0/tmp_reg[45]  ( .D(n1924), .CK(clk), .Q(ssrms0_out[45]) );
  DFFQX1TS \ssrms0/tmp_reg[43]  ( .D(n1922), .CK(clk), .Q(ssrms0_out[43]) );
  DFFQX1TS \ssrms0/tmp_reg[38]  ( .D(n1917), .CK(clk), .Q(ssrms0_out[38]) );
  DFFQX1TS \ssrms0/tmp_reg[36]  ( .D(n1915), .CK(clk), .Q(ssrms0_out[36]) );
  DFFQX1TS \ssrms0/tmp_reg[34]  ( .D(n1913), .CK(clk), .Q(ssrms0_out[34]) );
  DFFQX1TS \srmq/tmp_reg[59]  ( .D(n1778), .CK(clk), .Q(srmq_out[59]) );
  DFFQX1TS \srmq/tmp_reg[57]  ( .D(n1776), .CK(clk), .Q(srmq_out[57]) );
  DFFQX1TS \srmq/tmp_reg[55]  ( .D(n1774), .CK(clk), .Q(srmq_out[55]) );
  DFFQX1TS \srmq/tmp_reg[0]  ( .D(n1719), .CK(clk), .Q(srmq_out[0]) );
  DFFQX1TS \ssrms0/tmp_reg[35]  ( .D(n1914), .CK(clk), .Q(ssrms0_out[35]) );
  DFFQX1TS \srmq/tmp_reg[63]  ( .D(n1782), .CK(clk), .Q(srmq_out[63]) );
  DFFQX1TS \ssrms0/tmp_reg[37]  ( .D(n1916), .CK(clk), .Q(ssrms0_out[37]) );
  DFFQX1TS \srmq/tmp_reg[1]  ( .D(n1720), .CK(clk), .Q(srmq_out[1]) );
  DFFQX1TS \ssrms0/tmp_reg[42]  ( .D(n1921), .CK(clk), .Q(ssrms0_out[42]) );
  DFFQX1TS \ssrms0/tmp_reg[33]  ( .D(n1912), .CK(clk), .Q(ssrms0_out[33]) );
  DFFQX1TS \ssrms0/tmp_reg[39]  ( .D(n1918), .CK(clk), .Q(ssrms0_out[39]) );
  DFFQX1TS \ssrms0/tmp_reg[41]  ( .D(n1920), .CK(clk), .Q(ssrms0_out[41]) );
  DFFQX1TS \ssrms0/tmp_reg[32]  ( .D(n1911), .CK(clk), .Q(ssrms0_out[32]) );
  DFFQX1TS \srmq/tmp_reg[50]  ( .D(n1769), .CK(clk), .Q(srmq_out[50]) );
  DFFQX1TS \srmq/tmp_reg[19]  ( .D(n1738), .CK(clk), .Q(srmq_out[19]) );
  DFFQX1TS \srmq/tmp_reg[13]  ( .D(n1732), .CK(clk), .Q(srmq_out[13]) );
  DFFQX1TS \srmq/tmp_reg[7]  ( .D(n1726), .CK(clk), .Q(srmq_out[7]) );
  DFFQX1TS \srmq/tmp_reg[5]  ( .D(n1724), .CK(clk), .Q(srmq_out[5]) );
  DFFQX1TS \srmq/tmp_reg[3]  ( .D(n1722), .CK(clk), .Q(srmq_out[3]) );
  DFFQX1TS \ssrms0/tmp_reg[62]  ( .D(n1941), .CK(clk), .Q(ssrms0_out[62]) );
  DFFQX1TS \ssrms0/tmp_reg[58]  ( .D(n1937), .CK(clk), .Q(ssrms0_out[58]) );
  DFFQX1TS \ssrms0/tmp_reg[54]  ( .D(n1933), .CK(clk), .Q(ssrms0_out[54]) );
  DFFQX1TS \ssrms0/tmp_reg[46]  ( .D(n1925), .CK(clk), .Q(ssrms0_out[46]) );
  DFFQX1TS \srmq/tmp_reg[53]  ( .D(n1772), .CK(clk), .Q(srmq_out[53]) );
  DFFQX1TS \srmq/tmp_reg[52]  ( .D(n1771), .CK(clk), .Q(srmq_out[52]) );
  DFFQX1TS \srmq/tmp_reg[51]  ( .D(n1770), .CK(clk), .Q(srmq_out[51]) );
  DFFQX1TS \srmq/tmp_reg[48]  ( .D(n1767), .CK(clk), .Q(srmq_out[48]) );
  DFFQX1TS \srmq/tmp_reg[22]  ( .D(n1741), .CK(clk), .Q(srmq_out[22]) );
  DFFQX1TS \srmq/tmp_reg[20]  ( .D(n1739), .CK(clk), .Q(srmq_out[20]) );
  DFFQX1TS \srmq/tmp_reg[18]  ( .D(n1737), .CK(clk), .Q(srmq_out[18]) );
  DFFQX1TS \srmq/tmp_reg[16]  ( .D(n1735), .CK(clk), .Q(srmq_out[16]) );
  DFFQX1TS \srmq/tmp_reg[15]  ( .D(n1734), .CK(clk), .Q(srmq_out[15]) );
  DFFQX1TS \srmq/tmp_reg[14]  ( .D(n1733), .CK(clk), .Q(srmq_out[14]) );
  DFFQX1TS \srmq/tmp_reg[12]  ( .D(n1731), .CK(clk), .Q(srmq_out[12]) );
  DFFQX1TS \srmq/tmp_reg[10]  ( .D(n1729), .CK(clk), .Q(srmq_out[10]) );
  DFFQX1TS \srmq/tmp_reg[9]  ( .D(n1728), .CK(clk), .Q(srmq_out[9]) );
  DFFQX1TS \srmq/tmp_reg[8]  ( .D(n1727), .CK(clk), .Q(srmq_out[8]) );
  DFFQX1TS \ssrms0/tmp_reg[60]  ( .D(n1939), .CK(clk), .Q(ssrms0_out[60]) );
  DFFQX1TS \ssrms0/tmp_reg[48]  ( .D(n1927), .CK(clk), .Q(ssrms0_out[48]) );
  DFFQX1TS \srmq/tmp_reg[62]  ( .D(n1781), .CK(clk), .Q(srmq_out[62]) );
  DFFQX1TS \ssrms0/tmp_reg[50]  ( .D(n1929), .CK(clk), .Q(ssrms0_out[50]) );
  DFFQX1TS \ssrms0/tmp_reg[44]  ( .D(n1923), .CK(clk), .Q(ssrms0_out[44]) );
  DFFQX1TS \srmq/tmp_reg[60]  ( .D(n1779), .CK(clk), .Q(srmq_out[60]) );
  DFFQX1TS \srmq/tmp_reg[58]  ( .D(n1777), .CK(clk), .Q(srmq_out[58]) );
  DFFQX1TS \srmq/tmp_reg[56]  ( .D(n1775), .CK(clk), .Q(srmq_out[56]) );
  DFFQX1TS \srmq/tmp_reg[54]  ( .D(n1773), .CK(clk), .Q(srmq_out[54]) );
  DFFQX1TS \srmq/tmp_reg[49]  ( .D(n1768), .CK(clk), .Q(srmq_out[49]) );
  DFFQX1TS \srmq/tmp_reg[46]  ( .D(n1765), .CK(clk), .Q(srmq_out[46]) );
  DFFQX1TS \srmq/tmp_reg[21]  ( .D(n1740), .CK(clk), .Q(srmq_out[21]) );
  DFFQX1TS \srmq/tmp_reg[17]  ( .D(n1736), .CK(clk), .Q(srmq_out[17]) );
  DFFQX1TS \srmq/tmp_reg[11]  ( .D(n1730), .CK(clk), .Q(srmq_out[11]) );
  DFFQX1TS \srmq/tmp_reg[6]  ( .D(n1725), .CK(clk), .Q(srmq_out[6]) );
  DFFQX1TS \srmq/tmp_reg[4]  ( .D(n1723), .CK(clk), .Q(srmq_out[4]) );
  DFFQX1TS \srmq/tmp_reg[2]  ( .D(n1721), .CK(clk), .Q(srmq_out[2]) );
  DFFQX1TS \ssrms0/tmp_reg[56]  ( .D(n1935), .CK(clk), .Q(ssrms0_out[56]) );
  DFFQX1TS \ssrms0/tmp_reg[52]  ( .D(n1931), .CK(clk), .Q(ssrms0_out[52]) );
  DFFQX1TS \srmq/tmp_reg[45]  ( .D(n1764), .CK(clk), .Q(srmq_out[45]) );
  DFFQX1TS \srmq/tmp_reg[42]  ( .D(n1761), .CK(clk), .Q(srmq_out[42]) );
  DFFQX1TS \srmq/tmp_reg[38]  ( .D(n1757), .CK(clk), .Q(srmq_out[38]) );
  DFFQX1TS \srmq/tmp_reg[34]  ( .D(n1753), .CK(clk), .Q(srmq_out[34]) );
  DFFQX1TS \srmq/tmp_reg[32]  ( .D(n1751), .CK(clk), .Q(srmq_out[32]) );
  DFFQX1TS \srmq/tmp_reg[29]  ( .D(n1748), .CK(clk), .Q(srmq_out[29]) );
  DFFQX1TS \srmq/tmp_reg[25]  ( .D(n1744), .CK(clk), .Q(srmq_out[25]) );
  DFFQX1TS \srmq/tmp_reg[23]  ( .D(n1742), .CK(clk), .Q(srmq_out[23]) );
  DFFQX1TS \srmq/tmp_reg[43]  ( .D(n1762), .CK(clk), .Q(srmq_out[43]) );
  DFFQX1TS \srmq/tmp_reg[41]  ( .D(n1760), .CK(clk), .Q(srmq_out[41]) );
  DFFQX1TS \srmq/tmp_reg[39]  ( .D(n1758), .CK(clk), .Q(srmq_out[39]) );
  DFFQX1TS \srmq/tmp_reg[36]  ( .D(n1755), .CK(clk), .Q(srmq_out[36]) );
  DFFQX1TS \srmq/tmp_reg[35]  ( .D(n1754), .CK(clk), .Q(srmq_out[35]) );
  DFFQX1TS \srmq/tmp_reg[31]  ( .D(n1750), .CK(clk), .Q(srmq_out[31]) );
  DFFQX1TS \srmq/tmp_reg[27]  ( .D(n1746), .CK(clk), .Q(srmq_out[27]) );
  DFFQX1TS \srmq/tmp_reg[26]  ( .D(n1745), .CK(clk), .Q(srmq_out[26]) );
  DFFQX1TS \srmq/tmp_reg[44]  ( .D(n1763), .CK(clk), .Q(srmq_out[44]) );
  DFFQX1TS \srmq/tmp_reg[40]  ( .D(n1759), .CK(clk), .Q(srmq_out[40]) );
  DFFQX1TS \srmq/tmp_reg[37]  ( .D(n1756), .CK(clk), .Q(srmq_out[37]) );
  DFFQX1TS \srmq/tmp_reg[33]  ( .D(n1752), .CK(clk), .Q(srmq_out[33]) );
  DFFQX1TS \srmq/tmp_reg[30]  ( .D(n1749), .CK(clk), .Q(srmq_out[30]) );
  DFFQX1TS \srmq/tmp_reg[28]  ( .D(n1747), .CK(clk), .Q(srmq_out[28]) );
  DFFQX1TS \srmq/tmp_reg[24]  ( .D(n1743), .CK(clk), .Q(srmq_out[24]) );
  DFFQX1TS \ssrms0/tmp_reg[63]  ( .D(n1942), .CK(clk), .Q(ssrms0_out[63]) );
  DFFQX1TS \srmq/tmp_reg[47]  ( .D(n1766), .CK(clk), .Q(srmq_out[47]) );
  DFFQX1TS \count/data_out_reg[1]  ( .D(\count/N30 ), .CK(clk), .Q(
        count_out[1]) );
  DFFQX1TS \count/data_out_reg[0]  ( .D(\count/N29 ), .CK(clk), .Q(
        count_out[0]) );
  DFFQX1TS \regi/data_out_buffer_reg[1]  ( .D(n1685), .CK(clk), .Q(regi_out[1]) );
  DFFQX1TS \ssrms0/tmp_reg[31]  ( .D(n1910), .CK(clk), .Q(ssrms0_out[31]) );
  DFFQX1TS \ssrms0/tmp_reg[30]  ( .D(n1909), .CK(clk), .Q(ssrms0_out[30]) );
  DFFQX1TS \reges0/data_out_buffer_reg[31]  ( .D(n1649), .CK(clk), .Q(
        reges0_out[31]) );
  DFFQX1TS \reges0/data_out_buffer_reg[30]  ( .D(n1651), .CK(clk), .Q(
        reges0_out[30]) );
  DFFQX1TS \srres/tmp_reg[31]  ( .D(n1718), .CK(clk), .Q(regres_out[31]) );
  DFFQX1TS \reges0/data_out_buffer_reg[28]  ( .D(n1653), .CK(clk), .Q(
        reges0_out[28]) );
  DFFQX1TS \reges0/data_out_buffer_reg[29]  ( .D(n1652), .CK(clk), .Q(
        reges0_out[29]) );
  DFFQX1TS \ssrms0/tmp_reg[29]  ( .D(n1908), .CK(clk), .Q(ssrms0_out[29]) );
  DFFQX1TS \ssrms0/tmp_reg[28]  ( .D(n1907), .CK(clk), .Q(ssrms0_out[28]) );
  DFFQX1TS \srres/tmp_reg[28]  ( .D(n1715), .CK(clk), .Q(regres_out[28]) );
  DFFQX1TS \srres/tmp_reg[29]  ( .D(n1716), .CK(clk), .Q(regres_out[29]) );
  DFFQX1TS \srres/tmp_reg[30]  ( .D(n1717), .CK(clk), .Q(regres_out[30]) );
  DFFQX1TS \reges0/data_out_buffer_reg[27]  ( .D(n1654), .CK(clk), .Q(
        reges0_out[27]) );
  DFFQX1TS \reges0/data_out_buffer_reg[26]  ( .D(n1655), .CK(clk), .Q(
        reges0_out[26]) );
  DFFQX1TS \ssrms0/tmp_reg[27]  ( .D(n1906), .CK(clk), .Q(ssrms0_out[27]) );
  DFFQX1TS \ssrms0/tmp_reg[26]  ( .D(n1905), .CK(clk), .Q(ssrms0_out[26]) );
  DFFQX1TS \ssrms0/tmp_reg[25]  ( .D(n1904), .CK(clk), .Q(ssrms0_out[25]) );
  DFFQX1TS \srres/tmp_reg[27]  ( .D(n1714), .CK(clk), .Q(regres_out[27]) );
  DFFQX1TS \srres/tmp_reg[26]  ( .D(n1713), .CK(clk), .Q(regres_out[26]) );
  DFFQX1TS \reges0/data_out_buffer_reg[24]  ( .D(n1657), .CK(clk), .Q(
        reges0_out[24]) );
  DFFQX1TS \reges0/data_out_buffer_reg[25]  ( .D(n1656), .CK(clk), .Q(
        reges0_out[25]) );
  DFFQX1TS \srres/tmp_reg[24]  ( .D(n1711), .CK(clk), .Q(regres_out[24]) );
  DFFQX1TS \srres/tmp_reg[25]  ( .D(n1712), .CK(clk), .Q(regres_out[25]) );
  DFFQX1TS \ssrms0/tmp_reg[24]  ( .D(n1903), .CK(clk), .Q(ssrms0_out[24]) );
  DFFQX1TS \ssrms0/tmp_reg[23]  ( .D(n1902), .CK(clk), .Q(ssrms0_out[23]) );
  DFFQX1TS \ssrms0/tmp_reg[22]  ( .D(n1901), .CK(clk), .Q(ssrms0_out[22]) );
  DFFQX1TS \reges0/data_out_buffer_reg[20]  ( .D(n1661), .CK(clk), .Q(
        reges0_out[20]) );
  DFFQX1TS \reges0/data_out_buffer_reg[22]  ( .D(n1659), .CK(clk), .Q(
        reges0_out[22]) );
  DFFQX1TS \reges0/data_out_buffer_reg[23]  ( .D(n1658), .CK(clk), .Q(
        reges0_out[23]) );
  DFFQX1TS \srres/tmp_reg[23]  ( .D(n1710), .CK(clk), .Q(regres_out[23]) );
  DFFQX1TS \srres/tmp_reg[22]  ( .D(n1709), .CK(clk), .Q(regres_out[22]) );
  DFFQX1TS \ssrms0/tmp_reg[21]  ( .D(n1900), .CK(clk), .Q(ssrms0_out[21]) );
  DFFQX1TS \ssrms0/tmp_reg[20]  ( .D(n1899), .CK(clk), .Q(ssrms0_out[20]) );
  DFFQX1TS \reges0/data_out_buffer_reg[18]  ( .D(n1663), .CK(clk), .Q(
        reges0_out[18]) );
  DFFQX1TS \reges0/data_out_buffer_reg[19]  ( .D(n1662), .CK(clk), .Q(
        reges0_out[19]) );
  DFFQX1TS \reges0/data_out_buffer_reg[21]  ( .D(n1660), .CK(clk), .Q(
        reges0_out[21]) );
  DFFQX1TS \ssrms0/tmp_reg[18]  ( .D(n1897), .CK(clk), .Q(ssrms0_out[18]) );
  DFFQX1TS \srres/tmp_reg[19]  ( .D(n1706), .CK(clk), .Q(regres_out[19]) );
  DFFQX1TS \srres/tmp_reg[20]  ( .D(n1707), .CK(clk), .Q(regres_out[20]) );
  DFFQX1TS \srres/tmp_reg[18]  ( .D(n1705), .CK(clk), .Q(regres_out[18]) );
  DFFQX1TS \srres/tmp_reg[21]  ( .D(n1708), .CK(clk), .Q(regres_out[21]) );
  DFFQX1TS \ssrms0/tmp_reg[19]  ( .D(n1898), .CK(clk), .Q(ssrms0_out[19]) );
  DFFQX1TS \ssrms0/tmp_reg[17]  ( .D(n1896), .CK(clk), .Q(ssrms0_out[17]) );
  DFFQX1TS \reges0/data_out_buffer_reg[16]  ( .D(n1665), .CK(clk), .Q(
        reges0_out[16]) );
  DFFQX1TS \reges0/data_out_buffer_reg[17]  ( .D(n1664), .CK(clk), .Q(
        reges0_out[17]) );
  DFFQX1TS \srres/tmp_reg[16]  ( .D(n1703), .CK(clk), .Q(regres_out[16]) );
  DFFQX1TS \srres/tmp_reg[17]  ( .D(n1704), .CK(clk), .Q(regres_out[17]) );
  DFFQX1TS \ssrms0/tmp_reg[15]  ( .D(n1894), .CK(clk), .Q(ssrms0_out[15]) );
  DFFQX1TS \ssrms0/tmp_reg[14]  ( .D(n1893), .CK(clk), .Q(ssrms0_out[14]) );
  DFFQX1TS \ssrms0/tmp_reg[16]  ( .D(n1895), .CK(clk), .Q(ssrms0_out[16]) );
  DFFQX1TS \reges0/data_out_buffer_reg[13]  ( .D(n1668), .CK(clk), .Q(
        reges0_out[13]) );
  DFFQX1TS \reges0/data_out_buffer_reg[14]  ( .D(n1667), .CK(clk), .Q(
        reges0_out[14]) );
  DFFQX1TS \reges0/data_out_buffer_reg[15]  ( .D(n1666), .CK(clk), .Q(
        reges0_out[15]) );
  DFFQX1TS \srres/tmp_reg[15]  ( .D(n1702), .CK(clk), .Q(regres_out[15]) );
  DFFQX1TS \srres/tmp_reg[14]  ( .D(n1701), .CK(clk), .Q(regres_out[14]) );
  DFFQX1TS \ssrms0/tmp_reg[12]  ( .D(n1891), .CK(clk), .Q(ssrms0_out[12]) );
  DFFQX1TS \ssrms0/tmp_reg[13]  ( .D(n1892), .CK(clk), .Q(ssrms0_out[13]) );
  DFFQX1TS \reges0/data_out_buffer_reg[12]  ( .D(n1669), .CK(clk), .Q(
        reges0_out[12]) );
  DFFQX1TS \srres/tmp_reg[12]  ( .D(n1699), .CK(clk), .Q(regres_out[12]) );
  DFFQX1TS \srres/tmp_reg[13]  ( .D(n1700), .CK(clk), .Q(regres_out[13]) );
  DFFQX1TS \ssrms0/tmp_reg[11]  ( .D(n1890), .CK(clk), .Q(ssrms0_out[11]) );
  DFFQX1TS \ssrms0/tmp_reg[10]  ( .D(n1889), .CK(clk), .Q(ssrms0_out[10]) );
  DFFQX1TS \reges0/data_out_buffer_reg[8]  ( .D(n1673), .CK(clk), .Q(
        reges0_out[8]) );
  DFFQX1TS \reges0/data_out_buffer_reg[9]  ( .D(n1672), .CK(clk), .Q(
        reges0_out[9]) );
  DFFQX1TS \reges0/data_out_buffer_reg[10]  ( .D(n1671), .CK(clk), .Q(
        reges0_out[10]) );
  DFFQX1TS \reges0/data_out_buffer_reg[11]  ( .D(n1670), .CK(clk), .Q(
        reges0_out[11]) );
  DFFQX1TS \srres/tmp_reg[11]  ( .D(n1698), .CK(clk), .Q(regres_out[11]) );
  DFFQX1TS \srres/tmp_reg[10]  ( .D(n1697), .CK(clk), .Q(regres_out[10]) );
  DFFQX1TS \srres/tmp_reg[9]  ( .D(n1696), .CK(clk), .Q(regres_out[9]) );
  DFFQX1TS \ssrms0/tmp_reg[8]  ( .D(n1887), .CK(clk), .Q(ssrms0_out[8]) );
  DFFQX1TS \srres/tmp_reg[7]  ( .D(n1694), .CK(clk), .Q(regres_out[7]) );
  DFFQX1TS \reges0/data_out_buffer_reg[7]  ( .D(n1674), .CK(clk), .Q(
        reges0_out[7]) );
  DFFQX1TS \srres/tmp_reg[8]  ( .D(n1695), .CK(clk), .Q(regres_out[8]) );
  DFFQX1TS \ssrms0/tmp_reg[7]  ( .D(n1886), .CK(clk), .Q(ssrms0_out[7]) );
  DFFQX1TS \ssrms0/tmp_reg[6]  ( .D(n1885), .CK(clk), .Q(ssrms0_out[6]) );
  DFFQX1TS \reges0/data_out_buffer_reg[5]  ( .D(n1676), .CK(clk), .Q(
        reges0_out[5]) );
  DFFQX1TS \reges0/data_out_buffer_reg[6]  ( .D(n1675), .CK(clk), .Q(
        reges0_out[6]) );
  DFFQX1TS \srres/tmp_reg[6]  ( .D(n1693), .CK(clk), .Q(regres_out[6]) );
  DFFQX1TS \srres/tmp_reg[5]  ( .D(n1692), .CK(clk), .Q(regres_out[5]) );
  DFFQX1TS \ssrms0/tmp_reg[5]  ( .D(n1884), .CK(clk), .Q(ssrms0_out[5]) );
  DFFQX1TS \reges0/data_out_buffer_reg[4]  ( .D(n1677), .CK(clk), .Q(
        reges0_out[4]) );
  DFFQX1TS \srres/tmp_reg[4]  ( .D(n1691), .CK(clk), .Q(regres_out[4]) );
  DFFQX1TS \ssrms0/tmp_reg[3]  ( .D(n1882), .CK(clk), .Q(ssrms0_out[3]) );
  DFFQX1TS \ssrms0/tmp_reg[4]  ( .D(n1883), .CK(clk), .Q(ssrms0_out[4]) );
  DFFQX1TS \reges0/data_out_buffer_reg[3]  ( .D(n1678), .CK(clk), .Q(
        reges0_out[3]) );
  DFFQX1TS \srres/tmp_reg[2]  ( .D(n1689), .CK(clk), .Q(regres_out[2]) );
  DFFQX1TS \reges0/data_out_buffer_reg[2]  ( .D(n1679), .CK(clk), .Q(
        reges0_out[2]) );
  DFFQX1TS \ssrms0/tmp_reg[0]  ( .D(n1879), .CK(clk), .Q(ssrms0_out[0]) );
  DFFQX1TS \srres/tmp_reg[3]  ( .D(n1690), .CK(clk), .Q(regres_out[3]) );
  DFFQX1TS \ssrms0/tmp_reg[1]  ( .D(n1880), .CK(clk), .Q(ssrms0_out[1]) );
  DFFQX1TS \ssrms0/tmp_reg[2]  ( .D(n1881), .CK(clk), .Q(ssrms0_out[2]) );
  DFFQX1TS \srmt/tmp_reg[31]  ( .D(n1814), .CK(clk), .Q(srmt_out[31]) );
  DFFQX1TS \reges0/data_out_buffer_reg[0]  ( .D(n1681), .CK(clk), .Q(
        reges0_out[0]) );
  DFFQX1TS \reges0/data_out_buffer_reg[1]  ( .D(n1680), .CK(clk), .Q(
        reges0_out[1]) );
  DFFQX1TS \srres/tmp_reg[0]  ( .D(n1687), .CK(clk), .Q(regres_out[0]) );
  DFFQX1TS \srres/tmp_reg[1]  ( .D(n1688), .CK(clk), .Q(regres_out[1]) );
  DFFQX1TS \srmt/tmp_reg[29]  ( .D(n1812), .CK(clk), .Q(srmt_out[29]) );
  DFFQX1TS \srmt/tmp_reg[30]  ( .D(n1813), .CK(clk), .Q(srmt_out[30]) );
  DFFQX1TS \srmt/tmp_reg[27]  ( .D(n1810), .CK(clk), .Q(srmt_out[27]) );
  DFFQX1TS \srmt/tmp_reg[28]  ( .D(n1811), .CK(clk), .Q(srmt_out[28]) );
  DFFQX1TS \srmt/tmp_reg[25]  ( .D(n1808), .CK(clk), .Q(srmt_out[25]) );
  DFFQX1TS \srmt/tmp_reg[26]  ( .D(n1809), .CK(clk), .Q(srmt_out[26]) );
  DFFQX1TS \srmt/tmp_reg[23]  ( .D(n1806), .CK(clk), .Q(srmt_out[23]) );
  DFFQX1TS \srmt/tmp_reg[24]  ( .D(n1807), .CK(clk), .Q(srmt_out[24]) );
  DFFQX1TS \srmt/tmp_reg[21]  ( .D(n1804), .CK(clk), .Q(srmt_out[21]) );
  DFFQX1TS \srmt/tmp_reg[22]  ( .D(n1805), .CK(clk), .Q(srmt_out[22]) );
  DFFQX1TS \srmt/tmp_reg[19]  ( .D(n1802), .CK(clk), .Q(srmt_out[19]) );
  DFFQX1TS \srmt/tmp_reg[20]  ( .D(n1803), .CK(clk), .Q(srmt_out[20]) );
  DFFQX1TS \srmt/tmp_reg[18]  ( .D(n1801), .CK(clk), .Q(srmt_out[18]) );
  DFFQX1TS \srmt/tmp_reg[17]  ( .D(n1800), .CK(clk), .Q(srmt_out[17]) );
  DFFQX1TS \srmt/tmp_reg[16]  ( .D(n1799), .CK(clk), .Q(srmt_out[16]) );
  DFFQX1TS \srmt/tmp_reg[15]  ( .D(n1798), .CK(clk), .Q(srmt_out[15]) );
  DFFQX1TS \srmt/tmp_reg[14]  ( .D(n1797), .CK(clk), .Q(srmt_out[14]) );
  DFFQX1TS \srmt/tmp_reg[13]  ( .D(n1796), .CK(clk), .Q(srmt_out[13]) );
  DFFQX1TS \srmt/tmp_reg[12]  ( .D(n1795), .CK(clk), .Q(srmt_out[12]) );
  DFFQX1TS \srmt/tmp_reg[11]  ( .D(n1794), .CK(clk), .Q(srmt_out[11]) );
  DFFQX1TS \srmt/tmp_reg[10]  ( .D(n1793), .CK(clk), .Q(srmt_out[10]) );
  DFFQX1TS \srmt/tmp_reg[9]  ( .D(n1792), .CK(clk), .Q(srmt_out[9]) );
  DFFQX1TS \srmt/tmp_reg[8]  ( .D(n1791), .CK(clk), .Q(srmt_out[8]) );
  DFFQX1TS \srmt/tmp_reg[7]  ( .D(n1790), .CK(clk), .Q(srmt_out[7]) );
  DFFQX1TS \srmt/tmp_reg[6]  ( .D(n1789), .CK(clk), .Q(srmt_out[6]) );
  DFFQX1TS \srmt/tmp_reg[4]  ( .D(n1787), .CK(clk), .Q(srmt_out[4]) );
  DFFQX1TS \srmt/tmp_reg[5]  ( .D(n1788), .CK(clk), .Q(srmt_out[5]) );
  DFFQX1TS \srmt/tmp_reg[3]  ( .D(n1786), .CK(clk), .Q(srmt_out[3]) );
  DFFQX1TS \srmt/tmp_reg[2]  ( .D(n1785), .CK(clk), .Q(srmt_out[2]) );
  DFFQX1TS \srmt/tmp_reg[1]  ( .D(n1784), .CK(clk), .Q(srmt_out[1]) );
  DFFQX1TS \srmt/tmp_reg[0]  ( .D(n1783), .CK(clk), .Q(srmt_out[0]) );
  DFFXLTS \regi/data_out_buffer_reg[0]  ( .D(n1686), .CK(clk), .Q(regi_out[0]), 
        .QN(n4813) );
  EDFFX2TS \rege/data_out_buffer_reg[2]  ( .D(pe_out[2]), .E(reg_e), .CK(clk), 
        .Q(rege_out[2]), .QN(n4812) );
  EDFFX2TS \rege/data_out_buffer_reg[1]  ( .D(pe_out[1]), .E(reg_e), .CK(clk), 
        .Q(rege_out[1]), .QN(n4810) );
  EDFFX2TS \rege/data_out_buffer_reg[0]  ( .D(pe_out[0]), .E(reg_e), .CK(clk), 
        .Q(rege_out[0]), .QN(n4811) );
  EDFFX1TS \regsum/data_out_buffer_reg[7]  ( .D(m2_out[7]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[7]), .QN(n4793) );
  EDFFX1TS \regsum/data_out_buffer_reg[1]  ( .D(m2_out[1]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[1]), .QN(n4799) );
  EDFFX1TS \regsum/data_out_buffer_reg[20]  ( .D(m2_out[20]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[20]), .QN(n4795) );
  EDFFX1TS \regsum/data_out_buffer_reg[30]  ( .D(m2_out[30]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[30]), .QN(n4783) );
  EDFFX1TS \regsum/data_out_buffer_reg[11]  ( .D(m2_out[11]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[11]), .QN(n4792) );
  EDFFX1TS \regmb/data_out_buffer_reg[14]  ( .D(rf_bout[14]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[14]) );
  EDFFX1TS \regmb/data_out_buffer_reg[20]  ( .D(rf_bout[20]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[20]) );
  EDFFX1TS \rege/data_out_buffer_reg[3]  ( .D(pe_out[3]), .E(reg_e), .CK(clk), 
        .Q(rege_out[3]), .QN(n4772) );
  EDFFX1TS \rege/data_out_buffer_reg[4]  ( .D(pe_out[4]), .E(reg_e), .CK(clk), 
        .Q(rege_out[4]), .QN(n4778) );
  EDFFX1TS \reges/data_out_buffer_reg[0]  ( .D(regsum_out[23]), .E(reg_es), 
        .CK(clk), .Q(reges_out[0]), .QN(n4777) );
  EDFFX1TS \regindex/data_out_buffer_reg[5]  ( .D(m13_out[5]), .E(reg_index), 
        .CK(clk), .Q(regindex_out[5]), .QN(n4774) );
  EDFFX1TS \regindex/data_out_buffer_reg[4]  ( .D(m13_out[4]), .E(reg_index), 
        .CK(clk), .Q(regindex_out[4]), .QN(n4784) );
  EDFFX1TS \regsum/data_out_buffer_reg[26]  ( .D(m2_out[26]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[26]), .QN(n4782) );
  EDFFX1TS \regsum/data_out_buffer_reg[29]  ( .D(m2_out[29]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[29]), .QN(n4786) );
  EDFFX1TS \regsum/data_out_buffer_reg[25]  ( .D(m2_out[25]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[25]), .QN(n4781) );
  EDFFX1TS \regsum/data_out_buffer_reg[23]  ( .D(m2_out[23]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[23]), .QN(n4785) );
  EDFFX1TS \regsum/data_out_buffer_reg[24]  ( .D(m2_out[24]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[24]), .QN(n4775) );
  EDFFX1TS \regsum/data_out_buffer_reg[10]  ( .D(m2_out[10]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[10]), .QN(n4802) );
  EDFFX1TS \regsum/data_out_buffer_reg[3]  ( .D(m2_out[3]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[3]), .QN(n4794) );
  EDFFX1TS \regsum/data_out_buffer_reg[2]  ( .D(m2_out[2]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[2]), .QN(n4804) );
  EDFFX1TS \regsum/data_out_buffer_reg[0]  ( .D(m2_out[0]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[0]), .QN(n4789) );
  EDFFX1TS \regsum/data_out_buffer_reg[13]  ( .D(m2_out[13]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[13]), .QN(n4797) );
  EDFFX1TS \regsum/data_out_buffer_reg[22]  ( .D(m2_out[22]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[22]), .QN(n4790) );
  EDFFX1TS \regsum/data_out_buffer_reg[17]  ( .D(m2_out[17]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[17]), .QN(n4796) );
  EDFFX1TS \regsum/data_out_buffer_reg[15]  ( .D(m2_out[15]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[15]), .QN(n4791) );
  EDFFX1TS \regsum/data_out_buffer_reg[6]  ( .D(m2_out[6]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[6]), .QN(n4803) );
  EDFFX1TS \regsum/data_out_buffer_reg[5]  ( .D(m2_out[5]), .E(reg_sum), .CK(
        clk), .Q(regsum_out[5]), .QN(n4798) );
  EDFFX1TS \regsum/data_out_buffer_reg[28]  ( .D(m2_out[28]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[28]), .QN(n4776) );
  EDFFX1TS \regsum/data_out_buffer_reg[21]  ( .D(m2_out[21]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[21]), .QN(n4800) );
  EDFFX1TS \regsum/data_out_buffer_reg[18]  ( .D(m2_out[18]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[18]), .QN(n4801) );
  EDFFX1TS \regsum/data_out_buffer_reg[12]  ( .D(m2_out[12]), .E(reg_sum), 
        .CK(clk), .Q(regsum_out[12]), .QN(n4788) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[20]  ( .D(m3_out[20]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[20]), .QN(n4807) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[25]  ( .D(m3_out[25]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[25]), .QN(n4787) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[26]  ( .D(m3_out[26]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[26]), .QN(n4806) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[27]  ( .D(m3_out[27]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[27]), .QN(n4808) );
  EDFFX1TS \regcurrterm/data_out_buffer_reg[29]  ( .D(m3_out[29]), .E(
        reg_currterm), .CK(clk), .Q(regcurrterm_out[29]), .QN(n4805) );
  EDFFX1TS \regreg/data_out_buffer_reg[31]  ( .D(regsum_out[31]), .E(n1994), 
        .CK(clk), .Q(regreg_out[31]) );
  EDFFX1TS \regreg/data_out_buffer_reg[30]  ( .D(regsum_out[30]), .E(n1994), 
        .CK(clk), .Q(regreg_out[30]) );
  EDFFX1TS \regreg/data_out_buffer_reg[29]  ( .D(regsum_out[29]), .E(n1994), 
        .CK(clk), .Q(regreg_out[29]) );
  EDFFX1TS \regreg/data_out_buffer_reg[28]  ( .D(regsum_out[28]), .E(n1994), 
        .CK(clk), .Q(regreg_out[28]) );
  EDFFX1TS \regreg/data_out_buffer_reg[27]  ( .D(regsum_out[27]), .E(n1994), 
        .CK(clk), .Q(regreg_out[27]) );
  EDFFX1TS \regreg/data_out_buffer_reg[26]  ( .D(regsum_out[26]), .E(n1994), 
        .CK(clk), .Q(regreg_out[26]) );
  EDFFX1TS \regreg/data_out_buffer_reg[25]  ( .D(regsum_out[25]), .E(n1994), 
        .CK(clk), .Q(regreg_out[25]) );
  EDFFX1TS \regreg/data_out_buffer_reg[24]  ( .D(regsum_out[24]), .E(n1994), 
        .CK(clk), .Q(regreg_out[24]) );
  EDFFX1TS \regreg/data_out_buffer_reg[23]  ( .D(regsum_out[23]), .E(n1994), 
        .CK(clk), .Q(regreg_out[23]) );
  EDFFX1TS \regreg/data_out_buffer_reg[22]  ( .D(regsum_out[22]), .E(n1994), 
        .CK(clk), .Q(regreg_out[22]) );
  EDFFX1TS \regreg/data_out_buffer_reg[21]  ( .D(regsum_out[21]), .E(n1994), 
        .CK(clk), .Q(regreg_out[21]) );
  EDFFX1TS \regreg/data_out_buffer_reg[20]  ( .D(regsum_out[20]), .E(n1994), 
        .CK(clk), .Q(regreg_out[20]) );
  EDFFX1TS \regreg/data_out_buffer_reg[19]  ( .D(regsum_out[19]), .E(n1994), 
        .CK(clk), .Q(regreg_out[19]) );
  EDFFX1TS \regreg/data_out_buffer_reg[18]  ( .D(regsum_out[18]), .E(n1994), 
        .CK(clk), .Q(regreg_out[18]) );
  EDFFX1TS \regreg/data_out_buffer_reg[17]  ( .D(regsum_out[17]), .E(n1994), 
        .CK(clk), .Q(regreg_out[17]) );
  EDFFX1TS \regreg/data_out_buffer_reg[16]  ( .D(regsum_out[16]), .E(n1994), 
        .CK(clk), .Q(regreg_out[16]) );
  EDFFX1TS \regreg/data_out_buffer_reg[15]  ( .D(regsum_out[15]), .E(n1994), 
        .CK(clk), .Q(regreg_out[15]) );
  EDFFX1TS \regreg/data_out_buffer_reg[14]  ( .D(regsum_out[14]), .E(n1994), 
        .CK(clk), .Q(regreg_out[14]) );
  EDFFX1TS \regreg/data_out_buffer_reg[13]  ( .D(regsum_out[13]), .E(n1994), 
        .CK(clk), .Q(regreg_out[13]) );
  EDFFX1TS \regreg/data_out_buffer_reg[12]  ( .D(regsum_out[12]), .E(n1994), 
        .CK(clk), .Q(regreg_out[12]) );
  EDFFX1TS \regreg/data_out_buffer_reg[11]  ( .D(regsum_out[11]), .E(n1994), 
        .CK(clk), .Q(regreg_out[11]) );
  EDFFX1TS \regreg/data_out_buffer_reg[10]  ( .D(regsum_out[10]), .E(n1994), 
        .CK(clk), .Q(regreg_out[10]) );
  EDFFX1TS \regreg/data_out_buffer_reg[9]  ( .D(regsum_out[9]), .E(n1994), 
        .CK(clk), .Q(regreg_out[9]) );
  EDFFX1TS \regreg/data_out_buffer_reg[8]  ( .D(regsum_out[8]), .E(n1994), 
        .CK(clk), .Q(regreg_out[8]) );
  EDFFX1TS \regreg/data_out_buffer_reg[7]  ( .D(regsum_out[7]), .E(n1994), 
        .CK(clk), .Q(regreg_out[7]) );
  EDFFX1TS \regreg/data_out_buffer_reg[6]  ( .D(regsum_out[6]), .E(n1994), 
        .CK(clk), .Q(regreg_out[6]) );
  EDFFX1TS \regreg/data_out_buffer_reg[5]  ( .D(regsum_out[5]), .E(n1994), 
        .CK(clk), .Q(regreg_out[5]) );
  EDFFX1TS \regreg/data_out_buffer_reg[4]  ( .D(regsum_out[4]), .E(n1994), 
        .CK(clk), .Q(regreg_out[4]) );
  EDFFX1TS \regreg/data_out_buffer_reg[3]  ( .D(regsum_out[3]), .E(n1994), 
        .CK(clk), .Q(regreg_out[3]) );
  EDFFX1TS \regreg/data_out_buffer_reg[2]  ( .D(regsum_out[2]), .E(n1994), 
        .CK(clk), .Q(regreg_out[2]) );
  EDFFX1TS \regreg/data_out_buffer_reg[1]  ( .D(regsum_out[1]), .E(n1994), 
        .CK(clk), .Q(regreg_out[1]) );
  EDFFX1TS \regreg/data_out_buffer_reg[0]  ( .D(regsum_out[0]), .E(n1994), 
        .CK(clk), .Q(regreg_out[0]) );
  EDFFX1TS \regacc/data_out_buffer_reg[31]  ( .D(regsum_out[31]), .E(n1992), 
        .CK(clk), .Q(regacc_out[31]) );
  EDFFX1TS \regacc/data_out_buffer_reg[27]  ( .D(regsum_out[27]), .E(n1992), 
        .CK(clk), .Q(regacc_out[27]) );
  EDFFX1TS \regacc/data_out_buffer_reg[19]  ( .D(regsum_out[19]), .E(n1992), 
        .CK(clk), .Q(regacc_out[19]) );
  EDFFX1TS \regacc/data_out_buffer_reg[16]  ( .D(regsum_out[16]), .E(n1992), 
        .CK(clk), .Q(regacc_out[16]) );
  EDFFX1TS \regacc/data_out_buffer_reg[14]  ( .D(regsum_out[14]), .E(n1992), 
        .CK(clk), .Q(regacc_out[14]) );
  EDFFX1TS \regacc/data_out_buffer_reg[9]  ( .D(regsum_out[9]), .E(n1992), 
        .CK(clk), .Q(regacc_out[9]) );
  EDFFX1TS \regacc/data_out_buffer_reg[8]  ( .D(regsum_out[8]), .E(n1992), 
        .CK(clk), .Q(regacc_out[8]) );
  EDFFX1TS \regacc/data_out_buffer_reg[4]  ( .D(regsum_out[4]), .E(n1992), 
        .CK(clk), .Q(regacc_out[4]) );
  EDFFX1TS \regacc/data_out_buffer_reg[30]  ( .D(m1_out[30]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[30]) );
  EDFFX1TS \regacc/data_out_buffer_reg[29]  ( .D(m1_out[29]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[29]) );
  EDFFX1TS \regacc/data_out_buffer_reg[28]  ( .D(m1_out[28]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[28]) );
  EDFFX1TS \regacc/data_out_buffer_reg[26]  ( .D(m1_out[26]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[26]) );
  EDFFX1TS \regacc/data_out_buffer_reg[25]  ( .D(m1_out[25]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[25]) );
  EDFFX1TS \regacc/data_out_buffer_reg[24]  ( .D(m1_out[24]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[24]) );
  EDFFX1TS \regacc/data_out_buffer_reg[23]  ( .D(m1_out[23]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[23]) );
  EDFFX1TS \regacc/data_out_buffer_reg[22]  ( .D(m1_out[22]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[22]) );
  EDFFX1TS \regacc/data_out_buffer_reg[21]  ( .D(m1_out[21]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[21]) );
  EDFFX1TS \regacc/data_out_buffer_reg[20]  ( .D(m1_out[20]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[20]) );
  EDFFX1TS \regacc/data_out_buffer_reg[18]  ( .D(m1_out[18]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[18]) );
  EDFFX1TS \regacc/data_out_buffer_reg[17]  ( .D(m1_out[17]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[17]) );
  EDFFX1TS \regacc/data_out_buffer_reg[15]  ( .D(m1_out[15]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[15]) );
  EDFFX1TS \regacc/data_out_buffer_reg[13]  ( .D(m1_out[13]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[13]) );
  EDFFX1TS \regacc/data_out_buffer_reg[12]  ( .D(m1_out[12]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[12]) );
  EDFFX1TS \regacc/data_out_buffer_reg[11]  ( .D(m1_out[11]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[11]) );
  EDFFX1TS \regacc/data_out_buffer_reg[10]  ( .D(m1_out[10]), .E(reg_acc), 
        .CK(clk), .Q(regacc_out[10]) );
  EDFFX1TS \regacc/data_out_buffer_reg[7]  ( .D(m1_out[7]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[7]) );
  EDFFX1TS \regacc/data_out_buffer_reg[6]  ( .D(m1_out[6]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[6]) );
  EDFFX1TS \regacc/data_out_buffer_reg[5]  ( .D(m1_out[5]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[5]) );
  EDFFX1TS \regacc/data_out_buffer_reg[3]  ( .D(m1_out[3]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[3]) );
  EDFFX1TS \regacc/data_out_buffer_reg[2]  ( .D(m1_out[2]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[2]) );
  EDFFX1TS \regacc/data_out_buffer_reg[1]  ( .D(m1_out[1]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[1]) );
  EDFFX1TS \regacc/data_out_buffer_reg[0]  ( .D(m1_out[0]), .E(reg_acc), .CK(
        clk), .Q(regacc_out[0]) );
  EDFFX1TS \regst/data_out_buffer_reg  ( .D(regcurrterm_out[31]), .E(reg_st), 
        .CK(clk), .Q(regst_out) );
  EDFFX1TS \regss/data_out_buffer_reg  ( .D(regsum_out[31]), .E(reg_ss), .CK(
        clk), .Q(regss_out) );
  EDFFX1TS \regma/data_out_buffer_reg[22]  ( .D(rf_bout[22]), .E(reg_ma), .CK(
        clk), .Q(regma_out[22]) );
  EDFFX1TS \regma/data_out_buffer_reg[21]  ( .D(rf_bout[21]), .E(reg_ma), .CK(
        clk), .Q(regma_out[21]) );
  EDFFX1TS \regma/data_out_buffer_reg[20]  ( .D(rf_bout[20]), .E(reg_ma), .CK(
        clk), .Q(regma_out[20]) );
  EDFFX1TS \regma/data_out_buffer_reg[19]  ( .D(rf_bout[19]), .E(reg_ma), .CK(
        clk), .Q(regma_out[19]) );
  EDFFX1TS \regma/data_out_buffer_reg[18]  ( .D(rf_bout[18]), .E(reg_ma), .CK(
        clk), .Q(regma_out[18]) );
  EDFFX1TS \regma/data_out_buffer_reg[17]  ( .D(rf_bout[17]), .E(reg_ma), .CK(
        clk), .Q(regma_out[17]) );
  EDFFX1TS \regma/data_out_buffer_reg[16]  ( .D(rf_bout[16]), .E(reg_ma), .CK(
        clk), .Q(regma_out[16]) );
  EDFFX1TS \regma/data_out_buffer_reg[15]  ( .D(rf_bout[15]), .E(reg_ma), .CK(
        clk), .Q(regma_out[15]) );
  EDFFX1TS \regma/data_out_buffer_reg[14]  ( .D(rf_bout[14]), .E(reg_ma), .CK(
        clk), .Q(regma_out[14]) );
  EDFFX1TS \regma/data_out_buffer_reg[13]  ( .D(rf_bout[13]), .E(reg_ma), .CK(
        clk), .Q(regma_out[13]) );
  EDFFX1TS \regma/data_out_buffer_reg[12]  ( .D(rf_bout[12]), .E(reg_ma), .CK(
        clk), .Q(regma_out[12]) );
  EDFFX1TS \regma/data_out_buffer_reg[11]  ( .D(rf_bout[11]), .E(reg_ma), .CK(
        clk), .Q(regma_out[11]) );
  EDFFX1TS \regma/data_out_buffer_reg[10]  ( .D(rf_bout[10]), .E(reg_ma), .CK(
        clk), .Q(regma_out[10]) );
  EDFFX1TS \regma/data_out_buffer_reg[9]  ( .D(rf_bout[9]), .E(reg_ma), .CK(
        clk), .Q(regma_out[9]) );
  EDFFX1TS \regma/data_out_buffer_reg[8]  ( .D(rf_bout[8]), .E(reg_ma), .CK(
        clk), .Q(regma_out[8]) );
  EDFFX1TS \regma/data_out_buffer_reg[7]  ( .D(rf_bout[7]), .E(reg_ma), .CK(
        clk), .Q(regma_out[7]) );
  EDFFX1TS \regma/data_out_buffer_reg[6]  ( .D(rf_bout[6]), .E(reg_ma), .CK(
        clk), .Q(regma_out[6]) );
  EDFFX1TS \regma/data_out_buffer_reg[5]  ( .D(rf_bout[5]), .E(reg_ma), .CK(
        clk), .Q(regma_out[5]) );
  EDFFX1TS \regma/data_out_buffer_reg[4]  ( .D(rf_bout[4]), .E(reg_ma), .CK(
        clk), .Q(regma_out[4]) );
  EDFFX1TS \regma/data_out_buffer_reg[3]  ( .D(rf_bout[3]), .E(reg_ma), .CK(
        clk), .Q(regma_out[3]) );
  EDFFX1TS \regma/data_out_buffer_reg[2]  ( .D(rf_bout[2]), .E(reg_ma), .CK(
        clk), .Q(regma_out[2]) );
  EDFFX1TS \regma/data_out_buffer_reg[1]  ( .D(rf_bout[1]), .E(reg_ma), .CK(
        clk), .Q(regma_out[1]) );
  EDFFX1TS \regma/data_out_buffer_reg[0]  ( .D(rf_bout[0]), .E(reg_ma), .CK(
        clk), .Q(regma_out[0]) );
  EDFFX1TS \reget/data_out_buffer_reg[7]  ( .D(regcurrterm_out[30]), .E(reg_et), .CK(clk), .Q(reget_out[7]) );
  EDFFX1TS \reget/data_out_buffer_reg[6]  ( .D(regcurrterm_out[29]), .E(reg_et), .CK(clk), .Q(reget_out[6]) );
  EDFFX1TS \reget/data_out_buffer_reg[5]  ( .D(regcurrterm_out[28]), .E(reg_et), .CK(clk), .Q(reget_out[5]) );
  EDFFX1TS \reget/data_out_buffer_reg[4]  ( .D(regcurrterm_out[27]), .E(reg_et), .CK(clk), .Q(reget_out[4]) );
  EDFFX1TS \reget/data_out_buffer_reg[3]  ( .D(regcurrterm_out[26]), .E(reg_et), .CK(clk), .Q(reget_out[3]) );
  EDFFX1TS \reget/data_out_buffer_reg[2]  ( .D(regcurrterm_out[25]), .E(reg_et), .CK(clk), .Q(reget_out[2]) );
  EDFFX1TS \reget/data_out_buffer_reg[1]  ( .D(regcurrterm_out[24]), .E(reg_et), .CK(clk), .Q(reget_out[1]) );
  EDFFX1TS \reget/data_out_buffer_reg[0]  ( .D(regcurrterm_out[23]), .E(reg_et), .CK(clk), .Q(reget_out[0]) );
  EDFFX1TS \reges/data_out_buffer_reg[7]  ( .D(regsum_out[30]), .E(reg_es), 
        .CK(clk), .Q(reges_out[7]) );
  EDFFX1TS \reges/data_out_buffer_reg[6]  ( .D(regsum_out[29]), .E(reg_es), 
        .CK(clk), .Q(reges_out[6]) );
  EDFFX1TS \reges/data_out_buffer_reg[5]  ( .D(regsum_out[28]), .E(reg_es), 
        .CK(clk), .Q(reges_out[5]) );
  EDFFX1TS \reges/data_out_buffer_reg[4]  ( .D(regsum_out[27]), .E(reg_es), 
        .CK(clk), .Q(reges_out[4]) );
  EDFFX1TS \reges/data_out_buffer_reg[3]  ( .D(regsum_out[26]), .E(reg_es), 
        .CK(clk), .Q(reges_out[3]) );
  EDFFX1TS \reges/data_out_buffer_reg[2]  ( .D(regsum_out[25]), .E(reg_es), 
        .CK(clk), .Q(reges_out[2]) );
  EDFFX1TS \reges/data_out_buffer_reg[1]  ( .D(regsum_out[24]), .E(reg_es), 
        .CK(clk), .Q(reges_out[1]) );
  EDFFX1TS \regsa/data_out_buffer_reg  ( .D(rf_bout[31]), .E(reg_sa), .CK(clk), 
        .Q(regsa_out) );
  EDFFX1TS \regss0/data_out_buffer_reg  ( .D(\m6_out[0] ), .E(reg_ss0), .CK(
        clk), .Q(regss0_out) );
  EDFFX1TS \regea/data_out_buffer_reg[7]  ( .D(rf_bout[30]), .E(reg_ea), .CK(
        clk), .Q(regea_out[7]) );
  EDFFX1TS \regea/data_out_buffer_reg[6]  ( .D(rf_bout[29]), .E(reg_ea), .CK(
        clk), .Q(regea_out[6]) );
  EDFFX1TS \regea/data_out_buffer_reg[5]  ( .D(rf_bout[28]), .E(reg_ea), .CK(
        clk), .Q(regea_out[5]) );
  EDFFX1TS \regea/data_out_buffer_reg[4]  ( .D(rf_bout[27]), .E(reg_ea), .CK(
        clk), .Q(regea_out[4]) );
  EDFFX1TS \regea/data_out_buffer_reg[3]  ( .D(rf_bout[26]), .E(reg_ea), .CK(
        clk), .Q(regea_out[3]) );
  EDFFX1TS \regea/data_out_buffer_reg[2]  ( .D(rf_bout[25]), .E(reg_ea), .CK(
        clk), .Q(regea_out[2]) );
  EDFFX1TS \regea/data_out_buffer_reg[1]  ( .D(rf_bout[24]), .E(reg_ea), .CK(
        clk), .Q(regea_out[1]) );
  EDFFX1TS \regea/data_out_buffer_reg[0]  ( .D(rf_bout[23]), .E(reg_ea), .CK(
        clk), .Q(regea_out[0]) );
  EDFFX1TS \regmb/data_out_buffer_reg[22]  ( .D(rf_bout[22]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[22]) );
  EDFFX1TS \regmb/data_out_buffer_reg[21]  ( .D(rf_bout[21]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[21]) );
  EDFFX1TS \regmb/data_out_buffer_reg[19]  ( .D(rf_bout[19]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[19]) );
  EDFFX1TS \regmb/data_out_buffer_reg[18]  ( .D(rf_bout[18]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[18]) );
  EDFFX1TS \regmb/data_out_buffer_reg[17]  ( .D(rf_bout[17]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[17]) );
  EDFFX1TS \regmb/data_out_buffer_reg[16]  ( .D(rf_bout[16]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[16]) );
  EDFFX1TS \regmb/data_out_buffer_reg[15]  ( .D(rf_bout[15]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[15]) );
  EDFFX1TS \regmb/data_out_buffer_reg[13]  ( .D(rf_bout[13]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[13]) );
  EDFFX1TS \regmb/data_out_buffer_reg[12]  ( .D(rf_bout[12]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[12]) );
  EDFFX1TS \regmb/data_out_buffer_reg[11]  ( .D(rf_bout[11]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[11]) );
  EDFFX1TS \regmb/data_out_buffer_reg[10]  ( .D(rf_bout[10]), .E(reg_mb), .CK(
        clk), .Q(regmb_out[10]) );
  ADDFX1TS \DP_OP_117J3_124_765/U3  ( .A(n4819), .B(count_out[4]), .CI(
        \DP_OP_117J3_124_765/n3 ), .CO(\DP_OP_117J3_124_765/n2 ), .S(
        \C43/DATA3_4 ) );
  ADDFX1TS \DP_OP_117J3_124_765/U5  ( .A(n4819), .B(count_out[2]), .CI(
        \DP_OP_117J3_124_765/n5 ), .CO(\DP_OP_117J3_124_765/n4 ), .S(
        \C43/DATA3_2 ) );
  ADDFX1TS \DP_OP_117J3_124_765/U4  ( .A(n4819), .B(count_out[3]), .CI(
        \DP_OP_117J3_124_765/n4 ), .CO(\DP_OP_117J3_124_765/n3 ), .S(
        \C43/DATA3_3 ) );
  ADDFX1TS \DP_OP_117J3_124_765/U6  ( .A(n4819), .B(count_out[1]), .CI(
        count_out[0]), .CO(\DP_OP_117J3_124_765/n5 ), .S(\C43/DATA3_1 ) );
  NAND3X1TS U2333 ( .A(\alutwo/N324 ), .B(alu2[0]), .C(n2476), .Y(n4715) );
  NOR4XLTS U2334 ( .A(n2974), .B(n2597), .C(n2596), .D(n2595), .Y(n2949) );
  NOR2X2TS U2335 ( .A(n2398), .B(mux9[2]), .Y(n2630) );
  INVX1TS U2336 ( .A(n3076), .Y(n3073) );
  INVX1TS U2337 ( .A(n2981), .Y(n2978) );
  INVX1TS U2338 ( .A(n3019), .Y(n3016) );
  INVX1TS U2339 ( .A(n3058), .Y(n3055) );
  INVX1TS U2340 ( .A(n3037), .Y(n3034) );
  NOR2X4TS U2341 ( .A(mux17[2]), .B(n2436), .Y(n3104) );
  INVX3TS U2342 ( .A(n4117), .Y(n4274) );
  NOR3X2TS U2343 ( .A(\alutwo/N324 ), .B(alu2[1]), .C(alu2[0]), .Y(n2455) );
  OR2X2TS U2344 ( .A(n3880), .B(n3751), .Y(n4135) );
  NOR2X4TS U2345 ( .A(mux17[2]), .B(mux17[0]), .Y(n3106) );
  NOR2X2TS U2346 ( .A(n2403), .B(n2387), .Y(n2388) );
  INVX3TS U2347 ( .A(n3768), .Y(n4407) );
  AND3X2TS U2348 ( .A(\aluone/N324 ), .B(alu1[1]), .C(n3133), .Y(n2316) );
  INVX3TS U2349 ( .A(n3764), .Y(n4412) );
  INVX3TS U2350 ( .A(n4304), .Y(n1985) );
  CLKBUFX3TS U2351 ( .A(n4515), .Y(n4595) );
  INVX3TS U2352 ( .A(n3780), .Y(n4592) );
  NOR2BX2TS U2353 ( .AN(n4729), .B(n3174), .Y(n3175) );
  INVX3TS U2354 ( .A(n3788), .Y(n4597) );
  INVX3TS U2355 ( .A(n4484), .Y(n1987) );
  NOR2X4TS U2356 ( .A(counterii[1]), .B(n4417), .Y(n4473) );
  NOR2X4TS U2357 ( .A(n4418), .B(n4417), .Y(n4479) );
  NOR2X2TS U2358 ( .A(n1991), .B(mux14[0]), .Y(n3286) );
  NOR2X4TS U2359 ( .A(\sr_mt[0] ), .B(n4418), .Y(n4476) );
  NOR2X4TS U2360 ( .A(counterii[1]), .B(\sr_mt[0] ), .Y(n4483) );
  NOR2X4TS U2361 ( .A(sr_res[0]), .B(sr_res[1]), .Y(n4603) );
  INVX2TS U2362 ( .A(1'b1), .Y(rege_out[5]) );
  INVX2TS U2364 ( .A(1'b1), .Y(rege_out[6]) );
  INVX2TS U2366 ( .A(1'b1), .Y(rege_out[7]) );
  INVX2TS U2368 ( .A(1'b1), .Y(rege_out[8]) );
  INVX2TS U2370 ( .A(1'b1), .Y(rege_out[9]) );
  INVX2TS U2372 ( .A(1'b1), .Y(rege_out[10]) );
  INVX2TS U2374 ( .A(1'b1), .Y(rege_out[11]) );
  INVX2TS U2376 ( .A(1'b1), .Y(rege_out[12]) );
  INVX2TS U2378 ( .A(1'b1), .Y(rege_out[13]) );
  INVX2TS U2380 ( .A(1'b1), .Y(rege_out[14]) );
  INVX2TS U2382 ( .A(1'b1), .Y(rege_out[15]) );
  INVX2TS U2384 ( .A(1'b1), .Y(rege_out[16]) );
  INVX2TS U2386 ( .A(1'b1), .Y(rege_out[17]) );
  INVX2TS U2388 ( .A(1'b1), .Y(rege_out[18]) );
  INVX2TS U2390 ( .A(1'b1), .Y(rege_out[19]) );
  INVX2TS U2392 ( .A(1'b1), .Y(rege_out[20]) );
  INVX2TS U2394 ( .A(1'b1), .Y(rege_out[21]) );
  INVX2TS U2396 ( .A(1'b1), .Y(rege_out[22]) );
  INVX2TS U2398 ( .A(1'b1), .Y(rege_out[23]) );
  INVX2TS U2400 ( .A(1'b1), .Y(rege_out[24]) );
  INVX2TS U2402 ( .A(1'b1), .Y(rege_out[25]) );
  INVX2TS U2404 ( .A(1'b1), .Y(rege_out[26]) );
  INVX2TS U2406 ( .A(1'b1), .Y(rege_out[27]) );
  INVX2TS U2408 ( .A(1'b1), .Y(rege_out[28]) );
  INVX2TS U2410 ( .A(1'b1), .Y(rege_out[29]) );
  INVX2TS U2412 ( .A(1'b1), .Y(rege_out[30]) );
  INVX2TS U2414 ( .A(1'b1), .Y(rege_out[31]) );
  INVX2TS U2416 ( .A(1'b1), .Y(reget_out[8]) );
  INVX2TS U2418 ( .A(1'b1), .Y(reget_out[9]) );
  INVX2TS U2420 ( .A(1'b1), .Y(reget_out[10]) );
  INVX2TS U2422 ( .A(1'b1), .Y(reget_out[11]) );
  INVX2TS U2424 ( .A(1'b1), .Y(reget_out[12]) );
  INVX2TS U2426 ( .A(1'b1), .Y(reget_out[13]) );
  INVX2TS U2428 ( .A(1'b1), .Y(reget_out[14]) );
  INVX2TS U2430 ( .A(1'b1), .Y(reget_out[15]) );
  INVX2TS U2432 ( .A(1'b1), .Y(reget_out[16]) );
  INVX2TS U2434 ( .A(1'b1), .Y(reget_out[17]) );
  INVX2TS U2436 ( .A(1'b1), .Y(reget_out[18]) );
  INVX2TS U2438 ( .A(1'b1), .Y(reget_out[19]) );
  INVX2TS U2440 ( .A(1'b1), .Y(reget_out[20]) );
  INVX2TS U2442 ( .A(1'b1), .Y(reget_out[21]) );
  INVX2TS U2444 ( .A(1'b1), .Y(reget_out[22]) );
  INVX2TS U2446 ( .A(1'b1), .Y(reget_out[23]) );
  INVX2TS U2448 ( .A(1'b1), .Y(reget_out[24]) );
  INVX2TS U2450 ( .A(1'b1), .Y(reget_out[25]) );
  INVX2TS U2452 ( .A(1'b1), .Y(reget_out[26]) );
  INVX2TS U2454 ( .A(1'b1), .Y(reget_out[27]) );
  INVX2TS U2456 ( .A(1'b1), .Y(reget_out[28]) );
  INVX2TS U2458 ( .A(1'b1), .Y(reget_out[29]) );
  INVX2TS U2460 ( .A(1'b1), .Y(reget_out[30]) );
  INVX2TS U2462 ( .A(1'b1), .Y(reget_out[31]) );
  INVX2TS U2464 ( .A(1'b1), .Y(reges_out[8]) );
  INVX2TS U2466 ( .A(1'b1), .Y(reges_out[9]) );
  INVX2TS U2468 ( .A(1'b1), .Y(reges_out[10]) );
  INVX2TS U2470 ( .A(1'b1), .Y(reges_out[11]) );
  INVX2TS U2472 ( .A(1'b1), .Y(reges_out[12]) );
  INVX2TS U2474 ( .A(1'b1), .Y(reges_out[13]) );
  INVX2TS U2476 ( .A(1'b1), .Y(reges_out[14]) );
  INVX2TS U2478 ( .A(1'b1), .Y(reges_out[15]) );
  INVX2TS U2480 ( .A(1'b1), .Y(reges_out[16]) );
  INVX2TS U2482 ( .A(1'b1), .Y(reges_out[17]) );
  INVX2TS U2484 ( .A(1'b1), .Y(reges_out[18]) );
  INVX2TS U2486 ( .A(1'b1), .Y(reges_out[19]) );
  INVX2TS U2488 ( .A(1'b1), .Y(reges_out[20]) );
  INVX2TS U2490 ( .A(1'b1), .Y(reges_out[21]) );
  INVX2TS U2492 ( .A(1'b1), .Y(reges_out[22]) );
  INVX2TS U2494 ( .A(1'b1), .Y(reges_out[23]) );
  INVX2TS U2496 ( .A(1'b1), .Y(reges_out[24]) );
  INVX2TS U2498 ( .A(1'b1), .Y(reges_out[25]) );
  INVX2TS U2500 ( .A(1'b1), .Y(reges_out[26]) );
  INVX2TS U2502 ( .A(1'b1), .Y(reges_out[27]) );
  INVX2TS U2504 ( .A(1'b1), .Y(reges_out[28]) );
  INVX2TS U2506 ( .A(1'b1), .Y(reges_out[29]) );
  INVX2TS U2508 ( .A(1'b1), .Y(reges_out[30]) );
  INVX2TS U2510 ( .A(1'b1), .Y(reges_out[31]) );
  INVX2TS U2512 ( .A(1'b1), .Y(regi_out[2]) );
  INVX2TS U2514 ( .A(1'b1), .Y(regi_out[3]) );
  INVX2TS U2516 ( .A(1'b1), .Y(regi_out[4]) );
  INVX2TS U2518 ( .A(1'b1), .Y(regi_out[5]) );
  INVX2TS U2520 ( .A(1'b1), .Y(regeb_out[8]) );
  INVX2TS U2522 ( .A(1'b1), .Y(regeb_out[9]) );
  INVX2TS U2524 ( .A(1'b1), .Y(regeb_out[10]) );
  INVX2TS U2526 ( .A(1'b1), .Y(regeb_out[11]) );
  INVX2TS U2528 ( .A(1'b1), .Y(regeb_out[12]) );
  INVX2TS U2530 ( .A(1'b1), .Y(regeb_out[13]) );
  INVX2TS U2532 ( .A(1'b1), .Y(regeb_out[14]) );
  INVX2TS U2534 ( .A(1'b1), .Y(regeb_out[15]) );
  INVX2TS U2536 ( .A(1'b1), .Y(regeb_out[16]) );
  INVX2TS U2538 ( .A(1'b1), .Y(regeb_out[17]) );
  INVX2TS U2540 ( .A(1'b1), .Y(regeb_out[18]) );
  INVX2TS U2542 ( .A(1'b1), .Y(regeb_out[19]) );
  INVX2TS U2544 ( .A(1'b1), .Y(regeb_out[20]) );
  INVX2TS U2546 ( .A(1'b1), .Y(regeb_out[21]) );
  INVX2TS U2548 ( .A(1'b1), .Y(regeb_out[22]) );
  INVX2TS U2550 ( .A(1'b1), .Y(regeb_out[23]) );
  INVX2TS U2552 ( .A(1'b1), .Y(regeb_out[24]) );
  INVX2TS U2554 ( .A(1'b1), .Y(regeb_out[25]) );
  INVX2TS U2556 ( .A(1'b1), .Y(regeb_out[26]) );
  INVX2TS U2558 ( .A(1'b1), .Y(regeb_out[27]) );
  INVX2TS U2560 ( .A(1'b1), .Y(regeb_out[28]) );
  INVX2TS U2562 ( .A(1'b1), .Y(regeb_out[29]) );
  INVX2TS U2564 ( .A(1'b1), .Y(regeb_out[30]) );
  INVX2TS U2566 ( .A(1'b1), .Y(regeb_out[31]) );
  INVX2TS U2568 ( .A(1'b1), .Y(regec_out[8]) );
  INVX2TS U2570 ( .A(1'b1), .Y(regec_out[9]) );
  INVX2TS U2572 ( .A(1'b1), .Y(regec_out[10]) );
  INVX2TS U2574 ( .A(1'b1), .Y(regec_out[11]) );
  INVX2TS U2576 ( .A(1'b1), .Y(regec_out[12]) );
  INVX2TS U2578 ( .A(1'b1), .Y(regec_out[13]) );
  INVX2TS U2580 ( .A(1'b1), .Y(regec_out[14]) );
  INVX2TS U2582 ( .A(1'b1), .Y(regec_out[15]) );
  INVX2TS U2584 ( .A(1'b1), .Y(regec_out[16]) );
  INVX2TS U2586 ( .A(1'b1), .Y(regec_out[17]) );
  INVX2TS U2588 ( .A(1'b1), .Y(regec_out[18]) );
  INVX2TS U2590 ( .A(1'b1), .Y(regec_out[19]) );
  INVX2TS U2592 ( .A(1'b1), .Y(regec_out[20]) );
  INVX2TS U2594 ( .A(1'b1), .Y(regec_out[21]) );
  INVX2TS U2596 ( .A(1'b1), .Y(regec_out[22]) );
  INVX2TS U2598 ( .A(1'b1), .Y(regec_out[23]) );
  INVX2TS U2600 ( .A(1'b1), .Y(regec_out[24]) );
  INVX2TS U2602 ( .A(1'b1), .Y(regec_out[25]) );
  INVX2TS U2604 ( .A(1'b1), .Y(regec_out[26]) );
  INVX2TS U2606 ( .A(1'b1), .Y(regec_out[27]) );
  INVX2TS U2608 ( .A(1'b1), .Y(regec_out[28]) );
  INVX2TS U2610 ( .A(1'b1), .Y(regec_out[29]) );
  INVX2TS U2612 ( .A(1'b1), .Y(regec_out[30]) );
  INVX2TS U2614 ( .A(1'b1), .Y(regec_out[31]) );
  INVX2TS U2616 ( .A(1'b1), .Y(m18_out[8]) );
  INVX2TS U2618 ( .A(1'b1), .Y(m18_out[9]) );
  INVX2TS U2620 ( .A(1'b1), .Y(m18_out[10]) );
  INVX2TS U2622 ( .A(1'b1), .Y(m18_out[11]) );
  INVX2TS U2624 ( .A(1'b1), .Y(m18_out[12]) );
  INVX2TS U2626 ( .A(1'b1), .Y(m18_out[13]) );
  INVX2TS U2628 ( .A(1'b1), .Y(m18_out[14]) );
  INVX2TS U2630 ( .A(1'b1), .Y(m18_out[15]) );
  INVX2TS U2632 ( .A(1'b1), .Y(m18_out[16]) );
  INVX2TS U2634 ( .A(1'b1), .Y(m18_out[17]) );
  INVX2TS U2636 ( .A(1'b1), .Y(m18_out[18]) );
  INVX2TS U2638 ( .A(1'b1), .Y(m18_out[19]) );
  INVX2TS U2640 ( .A(1'b1), .Y(m18_out[20]) );
  INVX2TS U2642 ( .A(1'b1), .Y(m18_out[21]) );
  INVX2TS U2644 ( .A(1'b1), .Y(m18_out[22]) );
  INVX2TS U2646 ( .A(1'b1), .Y(m18_out[23]) );
  INVX2TS U2648 ( .A(1'b1), .Y(m18_out[24]) );
  INVX2TS U2650 ( .A(1'b1), .Y(m18_out[25]) );
  INVX2TS U2652 ( .A(1'b1), .Y(m18_out[26]) );
  INVX2TS U2654 ( .A(1'b1), .Y(m18_out[27]) );
  INVX2TS U2656 ( .A(1'b1), .Y(m18_out[28]) );
  INVX2TS U2658 ( .A(1'b1), .Y(m18_out[29]) );
  INVX2TS U2660 ( .A(1'b1), .Y(m18_out[30]) );
  INVX2TS U2662 ( .A(1'b1), .Y(m18_out[31]) );
  OAI21XLTS U2664 ( .A0(n2846), .A1(n2836), .B0(n2837), .Y(n2425) );
  OAI21XLTS U2665 ( .A0(n2422), .A1(n2421), .B0(n2420), .Y(n2423) );
  NOR2XLTS U2666 ( .A(n3094), .B(n3089), .Y(n3130) );
  NOR2XLTS U2667 ( .A(n3093), .B(n3103), .Y(n3135) );
  NOR2XLTS U2668 ( .A(n2758), .B(n2749), .Y(n2769) );
  NOR2XLTS U2669 ( .A(n2743), .B(n2753), .Y(n2763) );
  NOR2XLTS U2670 ( .A(n3069), .B(n2748), .Y(n3066) );
  NOR2XLTS U2671 ( .A(n2742), .B(n3079), .Y(n3068) );
  NOR2XLTS U2672 ( .A(n3051), .B(n2747), .Y(n3048) );
  NOR2XLTS U2673 ( .A(n2739), .B(n3061), .Y(n3050) );
  NAND2BXLTS U2674 ( .AN(n2683), .B(n2682), .Y(n2706) );
  OR2X1TS U2675 ( .A(n2659), .B(n2658), .Y(n2683) );
  NOR2XLTS U2676 ( .A(n3030), .B(n2642), .Y(n3027) );
  NOR2XLTS U2677 ( .A(n2636), .B(n3040), .Y(n3029) );
  NOR2XLTS U2678 ( .A(n2641), .B(n3012), .Y(n3009) );
  NOR2XLTS U2679 ( .A(n2633), .B(n3022), .Y(n3011) );
  NOR2XLTS U2680 ( .A(n2998), .B(n2612), .Y(n2952) );
  NOR2XLTS U2681 ( .A(n2603), .B(n2964), .Y(n2954) );
  NOR2XLTS U2682 ( .A(n2611), .B(n2974), .Y(n2971) );
  NOR2XLTS U2683 ( .A(n2600), .B(n2984), .Y(n2973) );
  NOR2XLTS U2684 ( .A(n2526), .B(n2525), .Y(n2527) );
  NOR2XLTS U2685 ( .A(n2509), .B(n2907), .Y(n2904) );
  NOR2XLTS U2686 ( .A(n2503), .B(n2917), .Y(n2906) );
  NOR2XLTS U2687 ( .A(n2508), .B(n2890), .Y(n2887) );
  NOR2XLTS U2688 ( .A(n2500), .B(n2900), .Y(n2889) );
  NOR2XLTS U2689 ( .A(n2858), .B(n2425), .Y(n2855) );
  NOR2XLTS U2690 ( .A(n2417), .B(n2868), .Y(n2857) );
  OAI21XLTS U2691 ( .A0(n3370), .A1(n3351), .B0(n3350), .Y(n2424) );
  NOR2XLTS U2692 ( .A(n3360), .B(n2423), .Y(n3351) );
  NOR2XLTS U2693 ( .A(n2826), .B(n2825), .Y(n2376) );
  OAI21XLTS U2694 ( .A0(n3622), .A1(n4660), .B0(n4722), .Y(n3683) );
  NOR2XLTS U2695 ( .A(n2469), .B(n3492), .Y(n3494) );
  NOR2XLTS U2696 ( .A(m17_out[4]), .B(n2472), .Y(n3452) );
  NOR2XLTS U2697 ( .A(n2464), .B(n3448), .Y(n3449) );
  NOR2XLTS U2698 ( .A(n2462), .B(n3330), .Y(n3331) );
  NOR2XLTS U2699 ( .A(n3129), .B(n3128), .Y(n3140) );
  NAND2BXLTS U2700 ( .AN(n3130), .B(n3131), .Y(n3095) );
  NAND2BXLTS U2701 ( .AN(n3135), .B(n3136), .Y(n3097) );
  NAND3XLTS U2702 ( .A(n2765), .B(n3064), .C(n2734), .Y(n2762) );
  NOR2XLTS U2703 ( .A(n2772), .B(n2782), .Y(n3088) );
  NOR2XLTS U2704 ( .A(n2768), .B(n2776), .Y(n3090) );
  NOR2XLTS U2705 ( .A(n2766), .B(n2765), .Y(n2767) );
  NAND2BXLTS U2706 ( .AN(n2763), .B(n2764), .Y(n2750) );
  NOR2XLTS U2707 ( .A(n2762), .B(n2735), .Y(n3082) );
  NOR2XLTS U2708 ( .A(n2740), .B(n3046), .Y(n2741) );
  NAND2BXLTS U2709 ( .AN(n3066), .B(n3065), .Y(n3070) );
  NAND2BXLTS U2710 ( .AN(n3068), .B(n3067), .Y(n3072) );
  NOR2XLTS U2711 ( .A(n2732), .B(n2731), .Y(n2734) );
  NAND4XLTS U2712 ( .A(n2949), .B(n2730), .C(n2729), .D(n3042), .Y(n2731) );
  NAND2BXLTS U2713 ( .AN(n3048), .B(n3047), .Y(n3052) );
  NAND2BXLTS U2714 ( .AN(n3050), .B(n3049), .Y(n3054) );
  NOR2XLTS U2715 ( .A(n3051), .B(n2728), .Y(n3042) );
  NOR2XLTS U2716 ( .A(n2706), .B(n2705), .Y(n2707) );
  NOR2XLTS U2717 ( .A(n2708), .B(n2716), .Y(n2737) );
  NOR2XLTS U2718 ( .A(n2712), .B(n2728), .Y(n2745) );
  NOR2XLTS U2719 ( .A(n2684), .B(n2692), .Y(n2703) );
  NOR2XLTS U2720 ( .A(n2688), .B(n2697), .Y(n2709) );
  XOR2XLTS U2721 ( .A(n2697), .B(n2706), .Y(n2692) );
  NOR2XLTS U2722 ( .A(n2732), .B(n3003), .Y(n3041) );
  NOR2XLTS U2723 ( .A(n2660), .B(n2668), .Y(n2680) );
  NOR2XLTS U2724 ( .A(n2682), .B(n2664), .Y(n2685) );
  XOR2XLTS U2725 ( .A(n2682), .B(n2683), .Y(n2668) );
  NOR2XLTS U2726 ( .A(n2637), .B(n2647), .Y(n2656) );
  NOR2XLTS U2727 ( .A(n2652), .B(n2643), .Y(n2662) );
  XOR2XLTS U2728 ( .A(n2652), .B(n2659), .Y(n2647) );
  NOR2XLTS U2729 ( .A(n2634), .B(n3007), .Y(n2635) );
  NAND2BXLTS U2730 ( .AN(n3027), .B(n3026), .Y(n3031) );
  NAND2BXLTS U2731 ( .AN(n3029), .B(n3028), .Y(n3033) );
  NOR2XLTS U2732 ( .A(n3012), .B(n2629), .Y(n2729) );
  NAND2BXLTS U2733 ( .AN(n3009), .B(n3008), .Y(n3013) );
  NAND2BXLTS U2734 ( .AN(n3011), .B(n3010), .Y(n3015) );
  NAND4XLTS U2735 ( .A(n2949), .B(n2730), .C(n2729), .D(n2948), .Y(n3003) );
  NOR2XLTS U2736 ( .A(n2607), .B(n2618), .Y(n2631) );
  NOR2XLTS U2737 ( .A(n2614), .B(n2629), .Y(n2638) );
  NOR2XLTS U2738 ( .A(n2604), .B(n2992), .Y(n2986) );
  NOR2XLTS U2739 ( .A(n2613), .B(n3001), .Y(n2987) );
  XOR2XLTS U2740 ( .A(n3001), .B(n2605), .Y(n2992) );
  NOR2XLTS U2741 ( .A(n3001), .B(n2998), .Y(n2730) );
  NOR2XLTS U2742 ( .A(n2601), .B(n2969), .Y(n2602) );
  NAND2BXLTS U2743 ( .AN(n2952), .B(n2951), .Y(n2955) );
  NAND2BXLTS U2744 ( .AN(n2954), .B(n2953), .Y(n2957) );
  NAND2BXLTS U2745 ( .AN(n2971), .B(n2970), .Y(n2975) );
  NAND2BXLTS U2746 ( .AN(n2973), .B(n2972), .Y(n2977) );
  NOR2XLTS U2747 ( .A(n2571), .B(n2570), .Y(n2572) );
  NOR2XLTS U2748 ( .A(n2573), .B(n2581), .Y(n2598) );
  NOR2XLTS U2749 ( .A(n2577), .B(n2597), .Y(n2608) );
  NOR2XLTS U2750 ( .A(n2551), .B(n2559), .Y(n2568) );
  NOR2XLTS U2751 ( .A(n2555), .B(n2564), .Y(n2574) );
  XOR2XLTS U2752 ( .A(n2564), .B(n2571), .Y(n2559) );
  NOR2XLTS U2753 ( .A(n2528), .B(n2536), .Y(n2549) );
  NOR2XLTS U2754 ( .A(n2532), .B(n2545), .Y(n2552) );
  OAI21XLTS U2755 ( .A0(n2527), .A1(n2545), .B0(n2571), .Y(n2536) );
  NOR2XLTS U2756 ( .A(n2504), .B(n2514), .Y(n2523) );
  NOR2XLTS U2757 ( .A(n2510), .B(n2519), .Y(n2529) );
  XOR2XLTS U2758 ( .A(n2519), .B(n2526), .Y(n2514) );
  NOR2XLTS U2759 ( .A(n2501), .B(n2885), .Y(n2502) );
  NAND2BXLTS U2760 ( .AN(n2904), .B(n2903), .Y(n2908) );
  NAND2BXLTS U2761 ( .AN(n2906), .B(n2905), .Y(n2910) );
  NAND2BXLTS U2762 ( .AN(n2499), .B(n2498), .Y(n2501) );
  NAND2BXLTS U2763 ( .AN(n2887), .B(n2886), .Y(n2891) );
  NAND2BXLTS U2764 ( .AN(n2889), .B(n2888), .Y(n2893) );
  NOR2XLTS U2765 ( .A(n2419), .B(n2430), .Y(n2496) );
  XOR2XLTS U2766 ( .A(n2498), .B(n2499), .Y(n2430) );
  NOR2XLTS U2767 ( .A(n3431), .B(n2426), .Y(n3417) );
  ADDFX1TS U2768 ( .A(n3432), .B(n3428), .CI(n3427), .CO(n2419), .S(n3429) );
  NOR2XLTS U2769 ( .A(n3407), .B(n3395), .Y(n2418) );
  NOR2XLTS U2770 ( .A(n3398), .B(n2415), .Y(n2389) );
  NOR2XLTS U2771 ( .A(n2858), .B(n2835), .Y(n2386) );
  NAND2BXLTS U2772 ( .AN(n2855), .B(n2854), .Y(n2859) );
  NAND2BXLTS U2773 ( .AN(n2857), .B(n2856), .Y(n2861) );
  NOR2XLTS U2774 ( .A(n2850), .B(n2413), .Y(n2416) );
  NOR2XLTS U2775 ( .A(n2835), .B(n2424), .Y(n2836) );
  NOR2XLTS U2776 ( .A(n2414), .B(n2849), .Y(n2838) );
  XOR2XLTS U2777 ( .A(n3352), .B(n3361), .Y(n3363) );
  NAND2BXLTS U2778 ( .AN(n3351), .B(n3350), .Y(n3362) );
  NAND3XLTS U2779 ( .A(n3366), .B(n3358), .C(n2376), .Y(n2833) );
  NOR2XLTS U2780 ( .A(n3358), .B(n2351), .Y(n2412) );
  ADDFX1TS U2781 ( .A(n2411), .B(n2410), .CI(n2422), .CO(n3352), .S(n2358) );
  AOI2BB1XLTS U2782 ( .A0N(n3357), .A1N(n2376), .B0(n3728), .Y(n3356) );
  OAI21XLTS U2783 ( .A0(n2352), .A1(n2826), .B0(n2351), .Y(n2814) );
  NOR2XLTS U2784 ( .A(n2818), .B(n2831), .Y(n2822) );
  NAND2BXLTS U2785 ( .AN(n2339), .B(n2338), .Y(n2324) );
  NOR2XLTS U2786 ( .A(n2327), .B(n3271), .Y(n2352) );
  NOR2XLTS U2787 ( .A(mux9[1]), .B(mux9[0]), .Y(n2401) );
  NOR3XLTS U2788 ( .A(mux9[1]), .B(mux8[2]), .C(n2298), .Y(n2702) );
  NOR3XLTS U2789 ( .A(mux9[1]), .B(mux8[2]), .C(mux8[0]), .Y(n2303) );
  NAND3XLTS U2790 ( .A(mux8[2]), .B(mux8[0]), .C(n2403), .Y(n2307) );
  NAND3XLTS U2791 ( .A(n3664), .B(n3645), .C(m17_out[28]), .Y(n3684) );
  NOR2XLTS U2792 ( .A(n3105), .B(n3112), .Y(n3118) );
  OAI21XLTS U2793 ( .A0(n3116), .A1(m17_out[27]), .B0(n3115), .Y(n3646) );
  NAND3XLTS U2794 ( .A(m17_out[24]), .B(m17_out[25]), .C(m17_out[26]), .Y(
        n3665) );
  NOR2XLTS U2795 ( .A(m17_out[22]), .B(n3609), .Y(n3622) );
  NOR2XLTS U2796 ( .A(n3665), .B(n3112), .Y(n3116) );
  NAND3XLTS U2797 ( .A(n3107), .B(m17_out[24]), .C(m17_out[25]), .Y(n3113) );
  AOI2BB1XLTS U2798 ( .A0N(n4715), .A1N(n3645), .B0(n3683), .Y(n3634) );
  NOR2XLTS U2799 ( .A(n3619), .B(n3109), .Y(n3111) );
  NOR2XLTS U2800 ( .A(m17_out[20]), .B(n3589), .Y(n3593) );
  NAND3XLTS U2801 ( .A(n3587), .B(m17_out[20]), .C(m17_out[21]), .Y(n3595) );
  OAI21XLTS U2802 ( .A0(n3110), .A1(m17_out[21]), .B0(n3109), .Y(n3596) );
  NOR2XLTS U2803 ( .A(n3608), .B(n3108), .Y(n3110) );
  NOR2XLTS U2804 ( .A(n3120), .B(n3119), .Y(n3587) );
  NOR2XLTS U2805 ( .A(m17_out[18]), .B(n3571), .Y(n2940) );
  NOR2XLTS U2806 ( .A(n3574), .B(n2932), .Y(n2934) );
  NAND3XLTS U2807 ( .A(n3541), .B(n4691), .C(n3539), .Y(n3571) );
  NOR2XLTS U2808 ( .A(n3541), .B(n2930), .Y(n2933) );
  NAND3XLTS U2809 ( .A(n3548), .B(m17_out[11]), .C(m17_out[12]), .Y(n3527) );
  NOR2XLTS U2810 ( .A(m17_out[15]), .B(n3565), .Y(n3539) );
  NAND4XLTS U2811 ( .A(n2929), .B(m17_out[13]), .C(m17_out[14]), .D(
        m17_out[15]), .Y(n2930) );
  NOR2XLTS U2812 ( .A(n3550), .B(n2919), .Y(n2931) );
  NOR2XLTS U2813 ( .A(m17_out[13]), .B(n4704), .Y(n3557) );
  NOR2XLTS U2814 ( .A(n3523), .B(n2938), .Y(n3547) );
  NOR2XLTS U2815 ( .A(m17_out[11]), .B(n3520), .Y(n3528) );
  NOR2XLTS U2816 ( .A(n2924), .B(n3486), .Y(n2927) );
  NOR2XLTS U2817 ( .A(m17_out[9]), .B(n4709), .Y(n3482) );
  OAI21XLTS U2818 ( .A0(n2925), .A1(m17_out[9]), .B0(n2924), .Y(n4712) );
  NOR2XLTS U2819 ( .A(m17_out[7]), .B(n2918), .Y(n3472) );
  NOR2XLTS U2820 ( .A(n2470), .B(n2484), .Y(n2923) );
  NOR2XLTS U2821 ( .A(n2920), .B(n4717), .Y(n2925) );
  NOR2XLTS U2822 ( .A(n2487), .B(n2475), .Y(n2936) );
  NAND2BXLTS U2823 ( .AN(n2923), .B(n2921), .Y(n2479) );
  AOI2BB2XLTS U2824 ( .B0(n3504), .B1(n3496), .A0N(n3496), .A1N(n3504), .Y(
        n3500) );
  NOR2XLTS U2825 ( .A(n2468), .B(n3504), .Y(n2467) );
  NOR2XLTS U2826 ( .A(n2473), .B(m17_out[5]), .Y(n3374) );
  NOR2XLTS U2827 ( .A(n2466), .B(n3385), .Y(n3375) );
  NAND3XLTS U2828 ( .A(n3456), .B(n3446), .C(n3445), .Y(n3378) );
  NAND2BXLTS U2829 ( .AN(n3452), .B(n3451), .Y(n3454) );
  NOR2XLTS U2830 ( .A(n2463), .B(n3456), .Y(n2465) );
  AOI2BB2XLTS U2831 ( .B0(n3333), .B1(m17_out[3]), .A0N(m17_out[3]), .A1N(
        n3333), .Y(n3335) );
  NOR2XLTS U2832 ( .A(n2460), .B(n3316), .Y(n3317) );
  OAI21XLTS U2833 ( .A0(n2869), .A1(n2471), .B0(n2870), .Y(n3320) );
  AND3X1TS U2834 ( .A(m17_out[2]), .B(m17_out[0]), .C(m17_out[1]), .Y(n2461)
         );
  NOR2XLTS U2835 ( .A(m17_out[0]), .B(m17_out[1]), .Y(n3309) );
  NOR2XLTS U2836 ( .A(n3303), .B(n2878), .Y(n2871) );
  NAND3XLTS U2837 ( .A(m18_out[0]), .B(m17_out[0]), .C(m17_out[1]), .Y(n2870)
         );
  NOR2XLTS U2838 ( .A(regeb_out[2]), .B(n2458), .Y(n3311) );
  XOR2XLTS U2839 ( .A(regss_out), .B(regst_out), .Y(xor3_out) );
  INVX2TS U2840 ( .A(reges0_out[5]), .Y(n3227) );
  INVX2TS U2841 ( .A(ssrms0_out[2]), .Y(n4286) );
  INVX2TS U2842 ( .A(ssrms0_out[5]), .Y(n4257) );
  INVX2TS U2843 ( .A(ssrms0_out[6]), .Y(n4248) );
  INVX2TS U2844 ( .A(regres_out[7]), .Y(n3442) );
  NOR2XLTS U2845 ( .A(n4663), .B(n3117), .Y(n3690) );
  ADDFX1TS U2846 ( .A(regi_out[1]), .B(regindex_out[1]), .CI(n3150), .CO(n3155), .S(n2809) );
  CLKAND2X2TS U2847 ( .A(regindex_out[0]), .B(regi_out[0]), .Y(n3150) );
  XOR2XLTS U2848 ( .A(n3735), .B(n3144), .Y(n3749) );
  NAND3XLTS U2849 ( .A(n3128), .B(n3085), .C(n3082), .Y(n3730) );
  OAI211XLTS U2850 ( .A0(n3740), .A1(n3739), .B0(n3738), .C0(n3737), .Y(n3745)
         );
  XOR2XLTS U2851 ( .A(n3094), .B(n3129), .Y(n3103) );
  OAI211XLTS U2852 ( .A0(n3739), .A1(n3097), .B0(n3096), .C0(n3737), .Y(n3099)
         );
  OAI21XLTS U2853 ( .A0(n3357), .A1(n3730), .B0(n3083), .Y(n3732) );
  NAND2BXLTS U2854 ( .AN(n3090), .B(n3091), .Y(n2773) );
  AOI211XLTS U2855 ( .A0(n3736), .A1(n2782), .B0(n3354), .C0(n2775), .Y(n2777)
         );
  OAI21XLTS U2856 ( .A0(n2767), .A1(n2782), .B0(n3129), .Y(n2776) );
  AOI211XLTS U2857 ( .A0(n3736), .A1(n2758), .B0(n3354), .C0(n2752), .Y(n2754)
         );
  XOR2XLTS U2858 ( .A(n2758), .B(n2766), .Y(n2753) );
  AO22XLTS U2859 ( .A0(n2750), .A1(n2316), .B0(n3419), .B1(n2751), .Y(n2756)
         );
  OAI211XLTS U2860 ( .A0(n3082), .A1(n2736), .B0(n3424), .C0(n3133), .Y(n2781)
         );
  OAI21XLTS U2861 ( .A0(n2741), .A1(n3069), .B0(n2766), .Y(n3079) );
  OAI211XLTS U2862 ( .A0(n3739), .A1(n3072), .B0(n3071), .C0(n3737), .Y(n3074)
         );
  OAI21XLTS U2863 ( .A0(n2734), .A1(n3357), .B0(n2733), .Y(n3062) );
  XOR2XLTS U2864 ( .A(n3051), .B(n2740), .Y(n3061) );
  OAI211XLTS U2865 ( .A0(n3739), .A1(n3054), .B0(n3053), .C0(n3737), .Y(n3056)
         );
  AOI211XLTS U2866 ( .A0(n3736), .A1(n2728), .B0(n3354), .C0(n2715), .Y(n2717)
         );
  OAI21XLTS U2867 ( .A0(n2707), .A1(n2728), .B0(n2740), .Y(n2716) );
  NAND2BXLTS U2868 ( .AN(n2737), .B(n2738), .Y(n2713) );
  NOR2XLTS U2869 ( .A(n2682), .B(n2678), .Y(n2679) );
  NAND2BXLTS U2870 ( .AN(n2703), .B(n2704), .Y(n2689) );
  AOI211XLTS U2871 ( .A0(n3736), .A1(n2697), .B0(n3354), .C0(n2691), .Y(n2693)
         );
  NOR2XLTS U2872 ( .A(n2947), .B(n3041), .Y(n2721) );
  NAND2BXLTS U2873 ( .AN(n2680), .B(n2681), .Y(n2665) );
  AOI211XLTS U2874 ( .A0(n3736), .A1(n2682), .B0(n3354), .C0(n2667), .Y(n2669)
         );
  NAND2BXLTS U2875 ( .AN(n2656), .B(n2657), .Y(n2644) );
  AOI211XLTS U2876 ( .A0(n3736), .A1(n2652), .B0(n3354), .C0(n2646), .Y(n2648)
         );
  AOI2BB1XLTS U2877 ( .A0N(n2678), .A1N(n3003), .B0(n2947), .Y(n2673) );
  OAI21XLTS U2878 ( .A0(n2635), .A1(n3030), .B0(n2659), .Y(n3040) );
  OAI211XLTS U2879 ( .A0(n3739), .A1(n3033), .B0(n3032), .C0(n3737), .Y(n3035)
         );
  OAI21XLTS U2880 ( .A0(n2729), .A1(n3357), .B0(n3004), .Y(n3023) );
  XOR2XLTS U2881 ( .A(n3012), .B(n2634), .Y(n3022) );
  OAI211XLTS U2882 ( .A0(n3739), .A1(n3015), .B0(n3014), .C0(n3737), .Y(n3017)
         );
  AOI2BB1XLTS U2883 ( .A0N(n3357), .A1N(n2730), .B0(n2997), .Y(n3004) );
  OAI21XLTS U2884 ( .A0(n2606), .A1(n2629), .B0(n2634), .Y(n2618) );
  AOI211XLTS U2885 ( .A0(n3736), .A1(n2629), .B0(n3354), .C0(n2617), .Y(n2619)
         );
  NAND2BXLTS U2886 ( .AN(n2631), .B(n2632), .Y(n2615) );
  NAND2BXLTS U2887 ( .AN(n2986), .B(n2985), .Y(n2989) );
  AOI211XLTS U2888 ( .A0(n3736), .A1(n3001), .B0(n3354), .C0(n2991), .Y(n2993)
         );
  AOI31XLTS U2889 ( .A0(n2730), .A1(n2949), .A2(n2948), .B0(n2947), .Y(n3002)
         );
  OAI21XLTS U2890 ( .A0(n2602), .A1(n2998), .B0(n2605), .Y(n2964) );
  OAI21XLTS U2891 ( .A0(n2949), .A1(n3357), .B0(n2733), .Y(n2997) );
  OAI211XLTS U2892 ( .A0(n3739), .A1(n2957), .B0(n2956), .C0(n3737), .Y(n2959)
         );
  XOR2XLTS U2893 ( .A(n2974), .B(n2601), .Y(n2984) );
  OAI211XLTS U2894 ( .A0(n3739), .A1(n2977), .B0(n2976), .C0(n3737), .Y(n2979)
         );
  AO21XLTS U2895 ( .A0(n2949), .A1(n2948), .B0(n2947), .Y(n2968) );
  OAI21XLTS U2896 ( .A0(n2572), .A1(n2597), .B0(n2601), .Y(n2581) );
  AOI211XLTS U2897 ( .A0(n3736), .A1(n2597), .B0(n3354), .C0(n2580), .Y(n2582)
         );
  NAND2BXLTS U2898 ( .AN(n2598), .B(n2599), .Y(n2578) );
  NAND2BXLTS U2899 ( .AN(n2568), .B(n2569), .Y(n2556) );
  AOI211XLTS U2900 ( .A0(n3736), .A1(n2564), .B0(n3354), .C0(n2558), .Y(n2560)
         );
  AOI31XLTS U2901 ( .A0(n2548), .A1(n2547), .A2(n2948), .B0(n2947), .Y(n2586)
         );
  NAND2BXLTS U2902 ( .AN(n2549), .B(n2550), .Y(n2533) );
  AOI211XLTS U2903 ( .A0(n3736), .A1(n2545), .B0(n3354), .C0(n2535), .Y(n2537)
         );
  NAND2BXLTS U2904 ( .AN(n2523), .B(n2524), .Y(n2511) );
  AOI211XLTS U2905 ( .A0(n3736), .A1(n2519), .B0(n3354), .C0(n2513), .Y(n2515)
         );
  OAI21XLTS U2906 ( .A0(n2502), .A1(n2907), .B0(n2526), .Y(n2917) );
  OAI211XLTS U2907 ( .A0(n3739), .A1(n2910), .B0(n2909), .C0(n3737), .Y(n2912)
         );
  XOR2XLTS U2908 ( .A(n2890), .B(n2501), .Y(n2900) );
  NOR3XLTS U2909 ( .A(n2498), .B(n2495), .C(n2494), .Y(n2883) );
  OAI211XLTS U2910 ( .A0(n3739), .A1(n2893), .B0(n2892), .C0(n3737), .Y(n2895)
         );
  NAND2BXLTS U2911 ( .AN(n2496), .B(n2497), .Y(n2427) );
  AOI211XLTS U2912 ( .A0(n3736), .A1(n2498), .B0(n3354), .C0(n2429), .Y(n2431)
         );
  OAI21XLTS U2913 ( .A0(n3421), .A1(n3427), .B0(n3419), .Y(n3420) );
  OAI21XLTS U2914 ( .A0(n2389), .A1(n3434), .B0(n2499), .Y(n3432) );
  OAI211XLTS U2915 ( .A0(n3739), .A1(n3401), .B0(n3400), .C0(n3737), .Y(n3402)
         );
  XOR2XLTS U2916 ( .A(n3395), .B(n3404), .Y(n3401) );
  OAI211XLTS U2917 ( .A0(n2371), .A1(n3442), .B0(n2370), .C0(n2369), .Y(n2372)
         );
  OAI211XLTS U2918 ( .A0(n2310), .A1(n2392), .B0(n2391), .C0(n2390), .Y(n3407)
         );
  INVX2TS U2919 ( .A(srmt_out[7]), .Y(n2392) );
  OAI21XLTS U2920 ( .A0(n2416), .A1(n2858), .B0(n2415), .Y(n2868) );
  OAI211XLTS U2921 ( .A0(n2398), .A1(n4248), .B0(n2394), .C0(n2393), .Y(n2395)
         );
  OAI211XLTS U2922 ( .A0(n3739), .A1(n2861), .B0(n2860), .C0(n3737), .Y(n2863)
         );
  NAND3XLTS U2923 ( .A(n2379), .B(n2378), .C(n2377), .Y(n2858) );
  AOI211XLTS U2924 ( .A0(\aluone/N324 ), .A1(n2495), .B0(alu1[1]), .C0(alu1[0]), .Y(n3397) );
  AO21XLTS U2925 ( .A0(n2850), .A1(n2413), .B0(n2416), .Y(n2849) );
  OAI211XLTS U2926 ( .A0(n2383), .A1(n3227), .B0(n2382), .C0(n2381), .Y(n2384)
         );
  AOI211XLTS U2927 ( .A0(n2316), .A1(n2842), .B0(n3354), .C0(n2840), .Y(n2841)
         );
  OAI211XLTS U2928 ( .A0(n2398), .A1(n4257), .B0(n2397), .C0(n2396), .Y(n2399)
         );
  OAI21XLTS U2929 ( .A0(n2834), .A1(n3357), .B0(n2882), .Y(n2851) );
  AO22XLTS U2930 ( .A0(n3362), .A1(n3419), .B0(n2316), .B1(n3363), .Y(n3353)
         );
  OAI21XLTS U2931 ( .A0(n3357), .A1(n2833), .B0(n3083), .Y(n3365) );
  NAND3XLTS U2932 ( .A(n2375), .B(n2374), .C(n2373), .Y(n3360) );
  OAI21XLTS U2933 ( .A0(n3358), .A1(n3357), .B0(n3356), .Y(n3359) );
  AOI211XLTS U2934 ( .A0(n2409), .A1(reges_out[4]), .B0(n2408), .C0(n2407), 
        .Y(n3370) );
  NOR2XLTS U2935 ( .A(n2346), .B(n2360), .Y(n2421) );
  AOI211XLTS U2936 ( .A0(n2409), .A1(reges_out[3]), .B0(n2350), .C0(n2349), 
        .Y(n2422) );
  OAI211XLTS U2937 ( .A0(n2383), .A1(n3169), .B0(n2333), .C0(n2332), .Y(n2334)
         );
  OAI21XLTS U2938 ( .A0(n2340), .A1(n2339), .B0(n2338), .Y(n2818) );
  XOR2XLTS U2939 ( .A(n2813), .B(n2814), .Y(n2819) );
  NOR2XLTS U2940 ( .A(n2826), .B(n3741), .Y(n2816) );
  NAND3XLTS U2941 ( .A(n2337), .B(n2336), .C(n2335), .Y(n2826) );
  AO22XLTS U2942 ( .A0(n2825), .A1(n3729), .B0(n2831), .B1(n3736), .Y(n2827)
         );
  NAND4XLTS U2943 ( .A(n2344), .B(n2343), .C(n2342), .D(n2341), .Y(n2831) );
  OAI211XLTS U2944 ( .A0(n2383), .A1(n2301), .B0(n2300), .C0(n2299), .Y(n2302)
         );
  NAND3XLTS U2945 ( .A(n3424), .B(n2736), .C(n3133), .Y(n3083) );
  AOI2BB1XLTS U2946 ( .A0N(n2403), .A1N(regms_out[1]), .B0(n2387), .Y(n2315)
         );
  OAI211XLTS U2947 ( .A0(n2406), .A1(n4810), .B0(n2313), .C0(n2312), .Y(n2314)
         );
  OAI211XLTS U2948 ( .A0(n2327), .A1(n3422), .B0(n2326), .C0(n3737), .Y(n2328)
         );
  NAND2BXLTS U2949 ( .AN(n2352), .B(n2825), .Y(n2355) );
  NOR2XLTS U2950 ( .A(n4811), .B(n2406), .Y(n2321) );
  OAI211XLTS U2951 ( .A0(n2319), .A1(n4777), .B0(n2318), .C0(n2317), .Y(n2320)
         );
  OAI21XLTS U2952 ( .A0(ssrms0_out[0]), .A1(mux9[2]), .B0(n2401), .Y(n2317) );
  NOR2XLTS U2953 ( .A(n2316), .B(n3419), .Y(n3266) );
  OAI211XLTS U2954 ( .A0(n2307), .A1(n2306), .B0(n2305), .C0(n2304), .Y(n2308)
         );
  INVX2TS U2955 ( .A(srmt_out[0]), .Y(n2306) );
  OAI21XLTS U2956 ( .A0(\aluone/N324 ), .A1(n3424), .B0(n3269), .Y(n3270) );
  AND3X1TS U2957 ( .A(alu1[1]), .B(\aluone/N324 ), .C(alu1[0]), .Y(n3403) );
  AOI2BB2XLTS U2958 ( .B0(n3690), .B1(m17_out[31]), .A0N(m17_out[31]), .A1N(
        n3690), .Y(n3691) );
  NOR2XLTS U2959 ( .A(n4663), .B(n4664), .Y(n3694) );
  NOR2XLTS U2960 ( .A(n4667), .B(n3676), .Y(n3692) );
  NOR2XLTS U2961 ( .A(n3639), .B(n3697), .Y(n3695) );
  NOR2XLTS U2962 ( .A(m17_out[29]), .B(n3686), .Y(n4661) );
  OAI21XLTS U2963 ( .A0(m17_out[29]), .A1(n4715), .B0(n3696), .Y(n4659) );
  OAI21XLTS U2964 ( .A0(n3118), .A1(m17_out[29]), .B0(n3117), .Y(n3677) );
  NOR2XLTS U2965 ( .A(n4715), .B(n3684), .Y(n3682) );
  NAND3XLTS U2966 ( .A(n3671), .B(n3670), .C(n4677), .Y(n3679) );
  NOR2XLTS U2967 ( .A(n3666), .B(n3665), .Y(n3664) );
  NOR2XLTS U2968 ( .A(m17_out[26]), .B(m17_out[27]), .Y(n3663) );
  NOR2XLTS U2969 ( .A(n3662), .B(n3661), .Y(n3678) );
  OAI21XLTS U2970 ( .A0(n3635), .A1(n4660), .B0(n3634), .Y(n3669) );
  OAI21XLTS U2971 ( .A0(n3647), .A1(n3646), .B0(n3661), .Y(n3651) );
  OAI21XLTS U2972 ( .A0(n3649), .A1(n4660), .B0(n3648), .Y(n3650) );
  NOR3XLTS U2973 ( .A(n3619), .B(n4676), .C(n3595), .Y(n3645) );
  NOR3XLTS U2974 ( .A(m17_out[26]), .B(m17_out[27]), .C(n3638), .Y(n3671) );
  NAND3XLTS U2975 ( .A(n4676), .B(n4679), .C(n3630), .Y(n3638) );
  NOR2XLTS U2976 ( .A(n3637), .B(n3636), .Y(n3647) );
  OAI21XLTS U2977 ( .A0(n3114), .A1(m17_out[25]), .B0(n3113), .Y(n3626) );
  NOR2XLTS U2978 ( .A(n4679), .B(n3112), .Y(n3114) );
  OAI21XLTS U2979 ( .A0(n4679), .A1(n4673), .B0(n4714), .Y(n3628) );
  NOR2XLTS U2980 ( .A(m17_out[23]), .B(m17_out[24]), .Y(n3627) );
  NOR2XLTS U2981 ( .A(n4672), .B(n4671), .Y(n4670) );
  OAI21XLTS U2982 ( .A0(n3111), .A1(m17_out[23]), .B0(n3112), .Y(n3620) );
  NOR2XLTS U2983 ( .A(n3606), .B(n3605), .Y(n3621) );
  NOR3XLTS U2984 ( .A(n3608), .B(n3611), .C(n3607), .Y(n3618) );
  OAI211XLTS U2985 ( .A0(n4660), .A1(n3609), .B0(n3619), .C0(n4714), .Y(n3617)
         );
  OAI21XLTS U2986 ( .A0(n3593), .A1(n4660), .B0(n4722), .Y(n3594) );
  OAI21XLTS U2987 ( .A0(n3597), .A1(n3596), .B0(n3605), .Y(n3598) );
  NOR2XLTS U2988 ( .A(n3584), .B(n3583), .Y(n3597) );
  NAND4XLTS U2989 ( .A(n4689), .B(n3585), .C(m17_out[19]), .D(m17_out[18]), 
        .Y(n3607) );
  NOR2XLTS U2990 ( .A(n2455), .B(m17_out[20]), .Y(n3586) );
  OAI211XLTS U2991 ( .A0(n3587), .A1(n4715), .B0(m17_out[20]), .C0(n4722), .Y(
        n3588) );
  OAI21XLTS U2992 ( .A0(n2940), .A1(n4660), .B0(n4722), .Y(n2941) );
  NAND3XLTS U2993 ( .A(n3585), .B(n4689), .C(m17_out[18]), .Y(n2943) );
  OAI21XLTS U2994 ( .A0(n2934), .A1(m17_out[19]), .B0(n3108), .Y(n2935) );
  NOR2XLTS U2995 ( .A(n4691), .B(n4686), .Y(n3585) );
  NOR2XLTS U2996 ( .A(n3570), .B(n4683), .Y(n3569) );
  OAI211XLTS U2997 ( .A0(n3585), .A1(n4715), .B0(n4722), .C0(n3572), .Y(n3573)
         );
  OAI21XLTS U2998 ( .A0(n2933), .A1(m17_out[17]), .B0(n2932), .Y(n4684) );
  OAI21XLTS U2999 ( .A0(n3571), .A1(n4660), .B0(n4714), .Y(n4687) );
  NOR2XLTS U3000 ( .A(n3538), .B(n3545), .Y(n4685) );
  NOR2XLTS U3001 ( .A(n3527), .B(n2939), .Y(n4688) );
  NAND3XLTS U3002 ( .A(m17_out[13]), .B(m17_out[14]), .C(m17_out[15]), .Y(
        n2939) );
  AO22XLTS U3003 ( .A0(n4689), .A1(n4688), .B0(n4710), .B1(n3539), .Y(n3542)
         );
  OAI21XLTS U3004 ( .A0(n2931), .A1(m17_out[15]), .B0(n2930), .Y(n3546) );
  NOR2XLTS U3005 ( .A(n3562), .B(n4697), .Y(n3561) );
  OAI21XLTS U3006 ( .A0(n3557), .A1(n4660), .B0(n3556), .Y(n3558) );
  NAND3XLTS U3007 ( .A(n4689), .B(n3548), .C(n3547), .Y(n4701) );
  OAI21XLTS U3008 ( .A0(n2929), .A1(m17_out[13]), .B0(n2928), .Y(n4698) );
  OAI21XLTS U3009 ( .A0(n3528), .A1(n4660), .B0(n3549), .Y(n3529) );
  NOR2XLTS U3010 ( .A(n4660), .B(n4704), .Y(n4700) );
  NOR2XLTS U3011 ( .A(n3486), .B(n3483), .Y(n3548) );
  NOR2XLTS U3012 ( .A(n3531), .B(n3530), .Y(n4699) );
  OAI21XLTS U3013 ( .A0(n2927), .A1(m17_out[11]), .B0(n2926), .Y(n3517) );
  NOR2XLTS U3014 ( .A(n3487), .B(n4711), .Y(n3518) );
  NOR2XLTS U3015 ( .A(n4717), .B(n4716), .Y(n4708) );
  NOR2XLTS U3016 ( .A(n4716), .B(n4715), .Y(n3474) );
  OAI211XLTS U3017 ( .A0(n3472), .A1(n4660), .B0(m17_out[8]), .C0(n4722), .Y(
        n3475) );
  NOR2XLTS U3018 ( .A(n3471), .B(n3470), .Y(n4713) );
  OAI211XLTS U3019 ( .A0(m18_out[7]), .A1(n2923), .B0(n2922), .C0(n2921), .Y(
        n3470) );
  NOR2XLTS U3020 ( .A(n4660), .B(n4709), .Y(n4718) );
  NOR2XLTS U3021 ( .A(m17_out[5]), .B(n3378), .Y(n3490) );
  OAI211XLTS U3022 ( .A0(n3504), .A1(n3503), .B0(n3502), .C0(n3501), .Y(n3505)
         );
  NOR2XLTS U3023 ( .A(regeb_out[6]), .B(n2458), .Y(n3507) );
  AOI2BB1XLTS U3024 ( .A0N(n2918), .A1N(n4660), .B0(n2455), .Y(n3510) );
  OAI211XLTS U3025 ( .A0(n3383), .A1(n3503), .B0(n3382), .C0(n3501), .Y(n3384)
         );
  NAND2BXLTS U3026 ( .AN(n3374), .B(n3373), .Y(n3381) );
  AOI31XLTS U3027 ( .A0(n4710), .A1(n3445), .A2(n3377), .B0(n2455), .Y(n3462)
         );
  NOR2XLTS U3028 ( .A(m17_out[4]), .B(m17_out[3]), .Y(n3377) );
  NOR2XLTS U3029 ( .A(regeb_out[4]), .B(n2458), .Y(n3459) );
  OAI211XLTS U3030 ( .A0(n3456), .A1(n3503), .B0(n3455), .C0(n3501), .Y(n3457)
         );
  NOR3XLTS U3031 ( .A(m17_out[2]), .B(m17_out[0]), .C(m17_out[1]), .Y(n3445)
         );
  NOR2XLTS U3032 ( .A(regeb_out[3]), .B(n2458), .Y(n3339) );
  OAI211XLTS U3033 ( .A0(n3446), .A1(n3503), .B0(n3336), .C0(n3501), .Y(n3337)
         );
  NAND2BXLTS U3034 ( .AN(n3320), .B(n4689), .Y(n3310) );
  OAI211XLTS U3035 ( .A0(n2876), .A1(n4715), .B0(n2875), .C0(n3501), .Y(n2877)
         );
  NOR2XLTS U3036 ( .A(m18_out[0]), .B(m17_out[0]), .Y(n3303) );
  NAND2BXLTS U3037 ( .AN(regeb_out[0]), .B(mux17[2]), .Y(m18_out[0]) );
  NOR2XLTS U3038 ( .A(n4774), .B(n3158), .Y(Coutadd) );
  OAI211XLTS U3039 ( .A0(n3749), .A1(n3748), .B0(n3747), .C0(n3746), .Y(
        aluone_out[31]) );
  MXI2XLTS U3040 ( .A(n3732), .B(n3731), .S0(n3735), .Y(n3747) );
  MXI2XLTS U3041 ( .A(n3745), .B(n3744), .S0(n3743), .Y(n3746) );
  AO21XLTS U3042 ( .A0(n3730), .A1(n3729), .B0(n3728), .Y(n3731) );
  OAI211XLTS U3043 ( .A0(n3103), .A1(n3748), .B0(n3102), .C0(n3101), .Y(
        aluone_out[30]) );
  OAI21XLTS U3044 ( .A0(n3085), .A1(n3357), .B0(n3084), .Y(n3086) );
  AO22XLTS U3045 ( .A0(n2773), .A1(n2316), .B0(n3419), .B1(n2774), .Y(n2779)
         );
  OAI211XLTS U3046 ( .A0(n3079), .A1(n3748), .B0(n3078), .C0(n3077), .Y(
        aluone_out[27]) );
  OAI211XLTS U3047 ( .A0(n3061), .A1(n3748), .B0(n3060), .C0(n3059), .Y(
        aluone_out[26]) );
  OAI21XLTS U3048 ( .A0(n3044), .A1(n3357), .B0(n3043), .Y(n3045) );
  AO22XLTS U3049 ( .A0(n2713), .A1(n2316), .B0(n3419), .B1(n2714), .Y(n2719)
         );
  AOI2BB1XLTS U3050 ( .A0N(n2679), .A1N(n3357), .B0(n3023), .Y(n2698) );
  AO22XLTS U3051 ( .A0(n2689), .A1(n2316), .B0(n3419), .B1(n2690), .Y(n2695)
         );
  AO22XLTS U3052 ( .A0(n2665), .A1(n2316), .B0(n3419), .B1(n2666), .Y(n2671)
         );
  AO22XLTS U3053 ( .A0(n2644), .A1(n2316), .B0(n3419), .B1(n2645), .Y(n2650)
         );
  OAI211XLTS U3054 ( .A0(n3040), .A1(n3748), .B0(n3039), .C0(n3038), .Y(
        aluone_out[21]) );
  OAI211XLTS U3055 ( .A0(n3022), .A1(n3748), .B0(n3021), .C0(n3020), .Y(
        aluone_out[20]) );
  OAI21XLTS U3056 ( .A0(n3005), .A1(n3357), .B0(n3004), .Y(n3006) );
  AO22XLTS U3057 ( .A0(n2615), .A1(n2316), .B0(n3419), .B1(n2616), .Y(n2621)
         );
  OAI211XLTS U3058 ( .A0(n3002), .A1(n3001), .B0(n3000), .C0(n2999), .Y(
        aluone_out[18]) );
  AO22XLTS U3059 ( .A0(n2989), .A1(n2316), .B0(n3419), .B1(n2990), .Y(n2995)
         );
  OAI211XLTS U3060 ( .A0(n2964), .A1(n3748), .B0(n2963), .C0(n2962), .Y(
        aluone_out[17]) );
  OAI211XLTS U3061 ( .A0(n2984), .A1(n3748), .B0(n2983), .C0(n2982), .Y(
        aluone_out[16]) );
  OAI21XLTS U3062 ( .A0(n2966), .A1(n3357), .B0(n2965), .Y(n2967) );
  AO22XLTS U3063 ( .A0(n2578), .A1(n2316), .B0(n3419), .B1(n2579), .Y(n2584)
         );
  AO22XLTS U3064 ( .A0(n2556), .A1(n2316), .B0(n3419), .B1(n2557), .Y(n2562)
         );
  AO22XLTS U3065 ( .A0(n2533), .A1(n2316), .B0(n3419), .B1(n2534), .Y(n2539)
         );
  AO22XLTS U3066 ( .A0(n2511), .A1(n2316), .B0(n3419), .B1(n2512), .Y(n2517)
         );
  OAI211XLTS U3067 ( .A0(n2917), .A1(n3748), .B0(n2916), .C0(n2915), .Y(
        aluone_out[11]) );
  OAI211XLTS U3068 ( .A0(n2900), .A1(n3748), .B0(n2899), .C0(n2898), .Y(
        aluone_out[10]) );
  OAI21XLTS U3069 ( .A0(n2883), .A1(n3357), .B0(n2882), .Y(n2884) );
  AO22XLTS U3070 ( .A0(n2427), .A1(n2316), .B0(n3419), .B1(n2428), .Y(n2433)
         );
  AOI211XLTS U3071 ( .A0(n3431), .A1(n3424), .B0(n3423), .C0(n3422), .Y(n3437)
         );
  OAI211XLTS U3072 ( .A0(n3408), .A1(n3407), .B0(n3406), .C0(n3405), .Y(
        aluone_out[7]) );
  AOI2BB2XLTS U3073 ( .B0(n2316), .B1(n3401), .A0N(n3741), .A1N(n3399), .Y(
        n3408) );
  OAI211XLTS U3074 ( .A0(n3748), .A1(n2868), .B0(n2867), .C0(n2866), .Y(
        aluone_out[6]) );
  NOR2XLTS U3075 ( .A(n2850), .B(n3357), .Y(n2852) );
  OAI211XLTS U3076 ( .A0(n3748), .A1(n2849), .B0(n2848), .C0(n2847), .Y(
        aluone_out[5]) );
  AOI31XLTS U3077 ( .A0(n2846), .A1(n3419), .A2(n2845), .B0(n2844), .Y(n2847)
         );
  OAI211XLTS U3078 ( .A0(n3370), .A1(n3369), .B0(n3368), .C0(n3367), .Y(
        aluone_out[4]) );
  AOI211XLTS U3079 ( .A0(n3355), .A1(n3360), .B0(n3354), .C0(n3353), .Y(n3369)
         );
  AOI31XLTS U3080 ( .A0(n2422), .A1(n3419), .A2(n2362), .B0(n2361), .Y(n2363)
         );
  OAI211XLTS U3081 ( .A0(n2832), .A1(n2831), .B0(n2830), .C0(n2829), .Y(
        aluone_out[2]) );
  OAI211XLTS U3082 ( .A0(n3748), .A1(n2355), .B0(n2331), .C0(n2330), .Y(
        aluone_out[1]) );
  OAI21XLTS U3083 ( .A0(n3275), .A1(n3737), .B0(n3274), .Y(aluone_out[0]) );
  OAI211XLTS U3084 ( .A0(n2456), .A1(n3701), .B0(n3700), .C0(n3699), .Y(
        alutwo_out[31]) );
  OAI21XLTS U3085 ( .A0(n4659), .A1(n3698), .B0(m17_out[31]), .Y(n3699) );
  AOI2BB1XLTS U3086 ( .A0N(n4661), .A1N(n4660), .B0(n4659), .Y(n4662) );
  OAI211XLTS U3087 ( .A0(n3689), .A1(n2456), .B0(n3688), .C0(n3687), .Y(
        alutwo_out[29]) );
  OAI211XLTS U3088 ( .A0(n3673), .A1(n2456), .B0(n3672), .C0(n3679), .Y(
        alutwo_out[28]) );
  OAI211XLTS U3089 ( .A0(n3654), .A1(m17_out[27]), .B0(n3653), .C0(n3652), .Y(
        alutwo_out[27]) );
  AOI31XLTS U3090 ( .A0(n3645), .A1(n4689), .A2(n3644), .B0(n2455), .Y(n3654)
         );
  OAI211XLTS U3091 ( .A0(n3649), .A1(n3648), .B0(n3643), .C0(n3642), .Y(
        alutwo_out[26]) );
  OAI21XLTS U3092 ( .A0(n2455), .A1(n3641), .B0(n3649), .Y(n3642) );
  OAI211XLTS U3093 ( .A0(n3633), .A1(n2456), .B0(n3632), .C0(n3631), .Y(
        alutwo_out[25]) );
  AOI211XLTS U3094 ( .A0(n4677), .A1(n4676), .B0(n4675), .C0(n4674), .Y(n4681)
         );
  AOI211XLTS U3095 ( .A0(n4710), .A1(m17_out[23]), .B0(n4679), .C0(n4678), .Y(
        n4680) );
  OAI21XLTS U3096 ( .A0(m17_out[23]), .A1(n3625), .B0(n3624), .Y(
        alutwo_out[23]) );
  OAI21XLTS U3097 ( .A0(n3621), .A1(n3620), .B0(n4671), .Y(n3623) );
  OAI21XLTS U3098 ( .A0(n3614), .A1(n2456), .B0(n3613), .Y(alutwo_out[22]) );
  OAI21XLTS U3099 ( .A0(n3618), .A1(n3617), .B0(n3612), .Y(n3613) );
  OAI211XLTS U3100 ( .A0(n3611), .A1(n4660), .B0(n3610), .C0(m17_out[22]), .Y(
        n3612) );
  OAI211XLTS U3101 ( .A0(n3611), .A1(n3610), .B0(n3601), .C0(n3600), .Y(
        alutwo_out[21]) );
  NAND2BXLTS U3102 ( .AN(n3609), .B(n4710), .Y(n3600) );
  OAI21XLTS U3103 ( .A0(n3608), .A1(n3607), .B0(n4714), .Y(n3599) );
  OAI21XLTS U3104 ( .A0(n3592), .A1(n2456), .B0(n3591), .Y(alutwo_out[20]) );
  OAI211XLTS U3105 ( .A0(n3589), .A1(n4660), .B0(n3586), .C0(n3607), .Y(n3590)
         );
  NOR2XLTS U3106 ( .A(n4660), .B(n3589), .Y(n2946) );
  OAI21XLTS U3107 ( .A0(n3577), .A1(n2456), .B0(n3576), .Y(alutwo_out[18]) );
  CLKAND2X2TS U3108 ( .A(n3585), .B(n4689), .Y(n3575) );
  AO21XLTS U3109 ( .A0(n4696), .A1(n4695), .B0(n4694), .Y(alutwo_out[17]) );
  OAI21XLTS U3110 ( .A0(n4685), .A1(n4684), .B0(n4683), .Y(n4695) );
  AOI31XLTS U3111 ( .A0(n4689), .A1(n4688), .A2(m17_out[16]), .B0(n4687), .Y(
        n4690) );
  OAI21XLTS U3112 ( .A0(n3544), .A1(n2456), .B0(n3543), .Y(alutwo_out[16]) );
  OAI21XLTS U3113 ( .A0(n4688), .A1(n4715), .B0(n4693), .Y(n3540) );
  OAI21XLTS U3114 ( .A0(n3555), .A1(n2456), .B0(n3554), .Y(alutwo_out[15]) );
  OAI211XLTS U3115 ( .A0(n3565), .A1(n4660), .B0(n3564), .C0(n3563), .Y(
        alutwo_out[14]) );
  OAI21XLTS U3116 ( .A0(n4703), .A1(n4701), .B0(n4714), .Y(n3559) );
  NOR4BXLTS U3117 ( .AN(n4701), .B(n2455), .C(n4700), .D(m17_out[13]), .Y(
        n4706) );
  AOI211XLTS U3118 ( .A0(n4710), .A1(n4704), .B0(n4703), .C0(n4702), .Y(n4705)
         );
  OAI211XLTS U3119 ( .A0(n3534), .A1(m17_out[12]), .B0(n3533), .C0(n3532), .Y(
        alutwo_out[12]) );
  AOI31XLTS U3120 ( .A0(n3548), .A1(n4689), .A2(m17_out[11]), .B0(n2455), .Y(
        n3534) );
  OAI21XLTS U3121 ( .A0(n3525), .A1(n2456), .B0(n3524), .Y(alutwo_out[11]) );
  OAI211XLTS U3122 ( .A0(n3520), .A1(n4660), .B0(n4714), .C0(n3519), .Y(n3521)
         );
  OAI211XLTS U3123 ( .A0(n3520), .A1(n4660), .B0(n3489), .C0(n3488), .Y(
        alutwo_out[10]) );
  OAI21XLTS U3124 ( .A0(n3483), .A1(n4715), .B0(n4714), .Y(n3484) );
  AOI2BB2XLTS U3125 ( .B0(n4710), .B1(n4709), .A0N(n4708), .A1N(n4715), .Y(
        n4724) );
  OAI211XLTS U3126 ( .A0(n3479), .A1(n2456), .B0(n3478), .C0(n3477), .Y(
        alutwo_out[8]) );
  OAI211XLTS U3127 ( .A0(n3510), .A1(m17_out[6]), .B0(n3509), .C0(n3508), .Y(
        alutwo_out[6]) );
  OAI21XLTS U3128 ( .A0(n3490), .A1(n4660), .B0(n4722), .Y(n3491) );
  OAI211XLTS U3129 ( .A0(n3388), .A1(m18_out[5]), .B0(n3387), .C0(n3386), .Y(
        alutwo_out[5]) );
  AO22XLTS U3130 ( .A0(n3383), .A1(n3462), .B0(m17_out[5]), .B1(n3379), .Y(
        n3387) );
  OAI211XLTS U3131 ( .A0(m17_out[4]), .A1(n3462), .B0(n3461), .C0(n3460), .Y(
        alutwo_out[4]) );
  OAI211XLTS U3132 ( .A0(n3342), .A1(m17_out[3]), .B0(n3341), .C0(n3340), .Y(
        alutwo_out[3]) );
  OAI21XLTS U3133 ( .A0(n3445), .A1(n4660), .B0(n4722), .Y(n3329) );
  OAI211XLTS U3134 ( .A0(n3326), .A1(n3325), .B0(n3324), .C0(n3323), .Y(
        alutwo_out[2]) );
  AOI211XLTS U3135 ( .A0(n4710), .A1(n3313), .B0(n3526), .C0(n3312), .Y(n3325)
         );
  OAI211XLTS U3136 ( .A0(n2881), .A1(m18_out[1]), .B0(n2880), .C0(n2879), .Y(
        alutwo_out[1]) );
  AOI2BB2XLTS U3137 ( .B0(n4689), .B1(n2876), .A0N(n3497), .A1N(n2874), .Y(
        n2881) );
  NOR3XLTS U3138 ( .A(alu1[1]), .B(n2736), .C(n3133), .Y(n2323) );
  OAI211XLTS U3139 ( .A0(n2406), .A1(n4772), .B0(n2348), .C0(n2347), .Y(n2349)
         );
  CLKBUFX2TS U3140 ( .A(n4821), .Y(regms_out[29]) );
  INVX2TS U3141 ( .A(n3403), .Y(n3748) );
  INVX2TS U3142 ( .A(mux9[1]), .Y(n2403) );
  NOR3X1TS U3143 ( .A(mux8[2]), .B(mux8[0]), .C(n2403), .Y(n2385) );
  INVX2TS U3144 ( .A(n2303), .Y(n2383) );
  INVX2TS U3145 ( .A(reges0_out[1]), .Y(n2301) );
  INVX2TS U3146 ( .A(n2307), .Y(n3125) );
  NOR4BX1TS U3147 ( .AN(mux8[2]), .B(\mux20[0] ), .C(mux9[1]), .D(mux8[0]), 
        .Y(n2699) );
  INVX2TS U3148 ( .A(n2699), .Y(n2371) );
  INVX2TS U3149 ( .A(n2371), .Y(n3122) );
  AOI22X1TS U3150 ( .A0(n3125), .A1(srmt_out[1]), .B0(n3122), .B1(
        regres_out[1]), .Y(n2300) );
  INVX2TS U3151 ( .A(mux8[0]), .Y(n2298) );
  NOR3X1TS U3152 ( .A(mux8[2]), .B(n2403), .C(n2298), .Y(n2380) );
  AOI22X1TS U3153 ( .A0(n2702), .A1(regms_out[1]), .B0(n2380), .B1(
        reges_out[1]), .Y(n2299) );
  AOI21X1TS U3154 ( .A0(n2385), .A1(reget_out[1]), .B0(n2302), .Y(n2327) );
  AOI22X1TS U3155 ( .A0(n3122), .A1(regres_out[0]), .B0(n2380), .B1(
        reges_out[0]), .Y(n2305) );
  AOI22X1TS U3156 ( .A0(n2303), .A1(reges0_out[0]), .B0(n2702), .B1(
        regms_out[0]), .Y(n2304) );
  AOI21X1TS U3157 ( .A0(n2385), .A1(reget_out[0]), .B0(n2308), .Y(n3271) );
  NAND2X1TS U3158 ( .A(n2327), .B(n3271), .Y(n2825) );
  INVX2TS U3159 ( .A(alu1[1]), .Y(n3424) );
  INVX2TS U3160 ( .A(alu1[0]), .Y(n3133) );
  NAND3X1TS U3161 ( .A(\aluone/N324 ), .B(n3424), .C(n3133), .Y(n3357) );
  INVX2TS U3162 ( .A(n3357), .Y(n3729) );
  INVX2TS U3163 ( .A(\aluone/N324 ), .Y(n2736) );
  NAND2X1TS U3164 ( .A(alu1[1]), .B(n2736), .Y(n2882) );
  INVX2TS U3165 ( .A(n2327), .Y(n2322) );
  AOI22X1TS U3166 ( .A0(n2327), .A1(n3083), .B0(n2882), .B1(n2322), .Y(n2309)
         );
  AOI21X1TS U3167 ( .A0(n3729), .A1(n2355), .B0(n2309), .Y(n2331) );
  INVX2TS U3168 ( .A(mux9[0]), .Y(n2311) );
  NAND2X1TS U3169 ( .A(n2311), .B(mux9[2]), .Y(n2387) );
  NAND2X1TS U3170 ( .A(mux9[2]), .B(n2403), .Y(n2406) );
  OR3X1TS U3171 ( .A(n2311), .B(mux9[1]), .C(mux9[2]), .Y(n2310) );
  INVX2TS U3172 ( .A(n2310), .Y(n3132) );
  NOR3X1TS U3173 ( .A(mux9[0]), .B(mux9[2]), .C(n2403), .Y(n2400) );
  AOI22X1TS U3174 ( .A0(n3132), .A1(srmt_out[1]), .B0(reget_out[1]), .B1(n2400), .Y(n2313) );
  NOR3X1TS U3175 ( .A(mux9[2]), .B(n2311), .C(n2403), .Y(n2409) );
  NAND2X1TS U3176 ( .A(reges_out[1]), .B(n2409), .Y(n2312) );
  AOI211XLTS U3177 ( .A0(n2401), .A1(ssrms0_out[1]), .B0(n2315), .C0(n2314), 
        .Y(n2340) );
  INVX2TS U3178 ( .A(n2316), .Y(n3739) );
  INVX2TS U3179 ( .A(n2387), .Y(n2402) );
  INVX2TS U3180 ( .A(n2409), .Y(n2319) );
  AOI22X1TS U3181 ( .A0(n3132), .A1(srmt_out[0]), .B0(reget_out[0]), .B1(n2400), .Y(n2318) );
  AOI211X1TS U3182 ( .A0(regms_out[0]), .A1(n2402), .B0(n2321), .C0(n2320), 
        .Y(n3267) );
  NAND2X1TS U3183 ( .A(n3271), .B(n3267), .Y(n2354) );
  INVX2TS U3184 ( .A(n2354), .Y(n3275) );
  AOI22X1TS U3185 ( .A0(n3275), .A1(n2322), .B0(n2355), .B1(n2354), .Y(n2325)
         );
  CLKBUFX2TS U3186 ( .A(n2323), .Y(n3419) );
  INVX2TS U3187 ( .A(n2323), .Y(n3741) );
  NAND2X1TS U3188 ( .A(n2327), .B(n3267), .Y(n2353) );
  NAND2X1TS U3189 ( .A(n2825), .B(n2353), .Y(n2339) );
  INVX2TS U3190 ( .A(n3267), .Y(n3268) );
  NAND2X1TS U3191 ( .A(n2352), .B(n3268), .Y(n2338) );
  OAI22X1TS U3192 ( .A0(n3739), .A1(n2325), .B0(n3741), .B1(n2324), .Y(n2329)
         );
  NOR2X1TS U3193 ( .A(\aluone/N324 ), .B(n3133), .Y(n3355) );
  INVX2TS U3194 ( .A(n3355), .Y(n3422) );
  AOI22X1TS U3195 ( .A0(n2316), .A1(n2325), .B0(n3419), .B1(n2324), .Y(n2326)
         );
  INVX2TS U3196 ( .A(n3422), .Y(n3736) );
  NAND2X1TS U3197 ( .A(alu1[1]), .B(n3736), .Y(n3737) );
  INVX2TS U3198 ( .A(n2340), .Y(n2356) );
  AOI22X1TS U3199 ( .A0(n2340), .A1(n2329), .B0(n2328), .B1(n2356), .Y(n2330)
         );
  INVX2TS U3200 ( .A(reges0_out[3]), .Y(n3169) );
  CLKBUFX2TS U3201 ( .A(n2702), .Y(n3123) );
  AOI22X1TS U3202 ( .A0(n3123), .A1(regms_out[3]), .B0(n3122), .B1(
        regres_out[3]), .Y(n2333) );
  AOI22X1TS U3203 ( .A0(n3125), .A1(srmt_out[3]), .B0(n2380), .B1(reges_out[3]), .Y(n2332) );
  AOI21X1TS U3204 ( .A0(n2385), .A1(reget_out[3]), .B0(n2334), .Y(n3358) );
  AOI22X1TS U3205 ( .A0(n3125), .A1(srmt_out[2]), .B0(n2380), .B1(reges_out[2]), .Y(n2337) );
  INVX2TS U3206 ( .A(n2383), .Y(n3124) );
  AOI22X1TS U3207 ( .A0(n3124), .A1(reges0_out[2]), .B0(n3123), .B1(
        regms_out[2]), .Y(n2336) );
  AOI22X1TS U3208 ( .A0(n3122), .A1(regres_out[2]), .B0(n2385), .B1(
        reget_out[2]), .Y(n2335) );
  INVX2TS U3209 ( .A(n2826), .Y(n2345) );
  INVX2TS U3210 ( .A(n2401), .Y(n2398) );
  OA22X1TS U3211 ( .A0(n4286), .A1(n2398), .B0(n4812), .B1(n2406), .Y(n2344)
         );
  AOI22X1TS U3212 ( .A0(reget_out[2]), .A1(n2400), .B0(reges_out[2]), .B1(
        n2409), .Y(n2343) );
  OAI21XLTS U3213 ( .A0(regms_out[2]), .A1(n2403), .B0(n2402), .Y(n2342) );
  NAND2X1TS U3214 ( .A(n3132), .B(srmt_out[2]), .Y(n2341) );
  NAND2X1TS U3215 ( .A(n2818), .B(n2831), .Y(n2823) );
  AOI21X1TS U3216 ( .A0(n2345), .A1(n2823), .B0(n2822), .Y(n2346) );
  INVX2TS U3217 ( .A(n3358), .Y(n2360) );
  NAND2X1TS U3218 ( .A(n2346), .B(n2360), .Y(n2420) );
  NOR2BX1TS U3219 ( .AN(n2420), .B(n2421), .Y(n2362) );
  OA22X1TS U3220 ( .A0(n3422), .A1(n3358), .B0(n3741), .B1(n2362), .Y(n2364)
         );
  NOR2BX1TS U3221 ( .AN(srmt_out[3]), .B(n2310), .Y(n2350) );
  AOI22X1TS U3222 ( .A0(ssrms0_out[3]), .A1(n2401), .B0(reget_out[3]), .B1(
        n2400), .Y(n2348) );
  OAI21XLTS U3223 ( .A0(regms_out[3]), .A1(n2403), .B0(n2402), .Y(n2347) );
  INVX2TS U3224 ( .A(n2882), .Y(n3728) );
  INVX2TS U3225 ( .A(n3083), .Y(n2947) );
  AOI21X1TS U3226 ( .A0(n3729), .A1(n2376), .B0(n2947), .Y(n2815) );
  NAND2X1TS U3227 ( .A(n2352), .B(n2826), .Y(n2351) );
  AOI21X1TS U3228 ( .A0(n3358), .A1(n2351), .B0(n2412), .Y(n2411) );
  AOI222XLTS U3229 ( .A0(n2356), .A1(n2355), .B0(n2356), .B1(n2354), .C0(n2355), .C1(n2353), .Y(n2813) );
  INVX2TS U3230 ( .A(n2813), .Y(n2357) );
  AOI222XLTS U3231 ( .A0(n2831), .A1(n2814), .B0(n2831), .B1(n2357), .C0(n2814), .C1(n2357), .Y(n2410) );
  AOI22X1TS U3232 ( .A0(n2316), .A1(n2358), .B0(n3403), .B1(n2411), .Y(n2359)
         );
  OAI221XLTS U3233 ( .A0(n3358), .A1(n3356), .B0(n2360), .B1(n2815), .C0(n2359), .Y(n2361) );
  AOI32X1TS U3234 ( .A0(n2364), .A1(n2363), .A2(n3737), .B0(n2422), .B1(n2363), 
        .Y(aluone_out[3]) );
  AOI22X1TS U3235 ( .A0(n3124), .A1(reges0_out[9]), .B0(n3123), .B1(
        regms_out[9]), .Y(n2365) );
  OAI2BB1X1TS U3236 ( .A0N(n3125), .A1N(srmt_out[9]), .B0(n2365), .Y(n2366) );
  AOI21X1TS U3237 ( .A0(n3122), .A1(regres_out[9]), .B0(n2366), .Y(n2507) );
  AOI22X1TS U3238 ( .A0(n3124), .A1(reges0_out[8]), .B0(n2699), .B1(
        regres_out[8]), .Y(n2368) );
  AOI22X1TS U3239 ( .A0(n3125), .A1(srmt_out[8]), .B0(n3123), .B1(regms_out[8]), .Y(n2367) );
  NAND2X1TS U3240 ( .A(n2368), .B(n2367), .Y(n3434) );
  INVX2TS U3241 ( .A(n3434), .Y(n3431) );
  AOI22X1TS U3242 ( .A0(n3125), .A1(srmt_out[7]), .B0(n2380), .B1(reges_out[7]), .Y(n2370) );
  AOI22X1TS U3243 ( .A0(n3123), .A1(regms_out[7]), .B0(n2385), .B1(
        reget_out[7]), .Y(n2369) );
  AOI21X1TS U3244 ( .A0(n3124), .A1(reges0_out[7]), .B0(n2372), .Y(n3398) );
  NAND2X1TS U3245 ( .A(n3431), .B(n3398), .Y(n2494) );
  AOI22X1TS U3246 ( .A0(n3123), .A1(regms_out[4]), .B0(n3122), .B1(
        regres_out[4]), .Y(n2375) );
  AOI22X1TS U3247 ( .A0(n3124), .A1(reges0_out[4]), .B0(n3125), .B1(
        srmt_out[4]), .Y(n2374) );
  AOI22X1TS U3248 ( .A0(n2380), .A1(reges_out[4]), .B0(n2385), .B1(
        reget_out[4]), .Y(n2373) );
  INVX2TS U3249 ( .A(n3360), .Y(n3366) );
  INVX2TS U3250 ( .A(n2833), .Y(n2834) );
  AOI22X1TS U3251 ( .A0(n2380), .A1(reges_out[6]), .B0(n2385), .B1(
        reget_out[6]), .Y(n2379) );
  AOI22X1TS U3252 ( .A0(n3124), .A1(reges0_out[6]), .B0(n3123), .B1(
        regms_out[6]), .Y(n2378) );
  AOI22X1TS U3253 ( .A0(n3125), .A1(srmt_out[6]), .B0(n3122), .B1(
        regres_out[6]), .Y(n2377) );
  AOI22X1TS U3254 ( .A0(n3122), .A1(regres_out[5]), .B0(n2380), .B1(
        reges_out[5]), .Y(n2382) );
  AOI22X1TS U3255 ( .A0(n3125), .A1(srmt_out[5]), .B0(n3123), .B1(regms_out[5]), .Y(n2381) );
  AOI21X1TS U3256 ( .A0(n2385), .A1(reget_out[5]), .B0(n2384), .Y(n2850) );
  INVX2TS U3257 ( .A(n2850), .Y(n2835) );
  AOI32X1TS U3258 ( .A0(n2834), .A1(n2882), .A2(n2386), .B0(n3357), .B1(n2882), 
        .Y(n3425) );
  AOI21X1TS U3259 ( .A0(n3729), .A1(n2494), .B0(n3425), .Y(n2435) );
  INVX2TS U3260 ( .A(n2507), .Y(n2498) );
  NAND2X1TS U3261 ( .A(n2386), .B(n2834), .Y(n2495) );
  OAI2BB1X1TS U3262 ( .A0N(n2494), .A1N(n3083), .B0(n3397), .Y(n3433) );
  AOI222X1TS U3263 ( .A0(ssrms0_out[9]), .A1(n2630), .B0(n2388), .B1(
        regms_out[9]), .C0(n3132), .C1(srmt_out[9]), .Y(n2506) );
  NAND2X1TS U3264 ( .A(n2412), .B(n3360), .Y(n2413) );
  NAND2X1TS U3265 ( .A(n2416), .B(n2858), .Y(n2415) );
  NAND2X1TS U3266 ( .A(n2389), .B(n3434), .Y(n2499) );
  AOI21X1TS U3267 ( .A0(n3398), .A1(n2415), .B0(n2389), .Y(n3404) );
  AOI22X1TS U3268 ( .A0(n2388), .A1(regms_out[7]), .B0(reget_out[7]), .B1(
        n2400), .Y(n2391) );
  AOI22X1TS U3269 ( .A0(ssrms0_out[7]), .A1(n2630), .B0(reges_out[7]), .B1(
        n2409), .Y(n2390) );
  AOI22X1TS U3270 ( .A0(reges_out[6]), .A1(n2409), .B0(reget_out[6]), .B1(
        n2400), .Y(n2394) );
  OAI21XLTS U3271 ( .A0(regms_out[6]), .A1(n2403), .B0(n2402), .Y(n2393) );
  AOI21X1TS U3272 ( .A0(n3132), .A1(srmt_out[6]), .B0(n2395), .Y(n2865) );
  AOI22X1TS U3273 ( .A0(n3132), .A1(srmt_out[5]), .B0(reget_out[5]), .B1(n2400), .Y(n2397) );
  OAI21XLTS U3274 ( .A0(regms_out[5]), .A1(n2403), .B0(n2402), .Y(n2396) );
  AOI21X1TS U3275 ( .A0(reges_out[5]), .A1(n2409), .B0(n2399), .Y(n2846) );
  NOR2BX1TS U3276 ( .AN(srmt_out[4]), .B(n2310), .Y(n2408) );
  AOI22X1TS U3277 ( .A0(ssrms0_out[4]), .A1(n2401), .B0(reget_out[4]), .B1(
        n2400), .Y(n2405) );
  OAI21XLTS U3278 ( .A0(regms_out[4]), .A1(n2403), .B0(n2402), .Y(n2404) );
  OAI211XLTS U3279 ( .A0(n2406), .A1(n4778), .B0(n2405), .C0(n2404), .Y(n2407)
         );
  OA21XLTS U3280 ( .A0(n2412), .A1(n3360), .B0(n2413), .Y(n3361) );
  AOI222XLTS U3281 ( .A0(n3370), .A1(n3352), .B0(n3370), .B1(n3361), .C0(n3352), .C1(n3361), .Y(n2414) );
  NAND2X1TS U3282 ( .A(n2414), .B(n2849), .Y(n2839) );
  AOI21X1TS U3283 ( .A0(n2846), .A1(n2839), .B0(n2838), .Y(n2417) );
  NAND2X1TS U3284 ( .A(n2417), .B(n2868), .Y(n2856) );
  AOI21X1TS U3285 ( .A0(n2865), .A1(n2856), .B0(n2857), .Y(n3395) );
  OAI2BB2XLTS U3286 ( .B0(n3404), .B1(n2418), .A0N(n3407), .A1N(n3395), .Y(
        n3428) );
  AOI222XLTS U3287 ( .A0(regms_out[8]), .A1(n2388), .B0(n2630), .B1(
        ssrms0_out[8]), .C0(srmt_out[8]), .C1(n3132), .Y(n3423) );
  INVX2TS U3288 ( .A(n3423), .Y(n3427) );
  NAND2X1TS U3289 ( .A(n2419), .B(n2430), .Y(n2497) );
  NAND2X1TS U3290 ( .A(n3360), .B(n2423), .Y(n3350) );
  NAND2X1TS U3291 ( .A(n2835), .B(n2424), .Y(n2837) );
  NAND2X1TS U3292 ( .A(n2858), .B(n2425), .Y(n2854) );
  AOI21X1TS U3293 ( .A0(n2865), .A1(n2854), .B0(n2855), .Y(n3396) );
  INVX2TS U3294 ( .A(n3398), .Y(n3426) );
  AOI222XLTS U3295 ( .A0(n3396), .A1(n3426), .B0(n3396), .B1(n3407), .C0(n3426), .C1(n3407), .Y(n2426) );
  NAND2X1TS U3296 ( .A(n3431), .B(n2426), .Y(n3418) );
  AOI21X1TS U3297 ( .A0(n3427), .A1(n3418), .B0(n3417), .Y(n2505) );
  OAI2BB2XLTS U3298 ( .B0(n2498), .B1(n2505), .A0N(n2505), .A1N(n2498), .Y(
        n2428) );
  INVX2TS U3299 ( .A(n3737), .Y(n3354) );
  OAI22X1TS U3300 ( .A0(n2428), .A1(n3741), .B0(n3739), .B1(n2427), .Y(n2429)
         );
  OAI22X1TS U3301 ( .A0(n2506), .A1(n2431), .B0(n2430), .B1(n3748), .Y(n2432)
         );
  AOI21X1TS U3302 ( .A0(n2506), .A1(n2433), .B0(n2432), .Y(n2434) );
  OAI221XLTS U3303 ( .A0(n2507), .A1(n2435), .B0(n2498), .B1(n3433), .C0(n2434), .Y(aluone_out[9]) );
  INVX2TS U3304 ( .A(mux17[2]), .Y(n2458) );
  NOR2X1TS U3305 ( .A(mux17[0]), .B(n2458), .Y(n2451) );
  INVX2TS U3306 ( .A(mux17[0]), .Y(n2436) );
  NOR2X1TS U3307 ( .A(n2458), .B(n2436), .Y(n2452) );
  AOI22X1TS U3308 ( .A0(n2451), .A1(regea_out[7]), .B0(regec_out[7]), .B1(
        n2452), .Y(n2438) );
  AOI22X1TS U3309 ( .A0(n3104), .A1(regep_out[7]), .B0(n3106), .B1(
        regeq_out[7]), .Y(n2437) );
  NAND2X1TS U3310 ( .A(n2438), .B(n2437), .Y(m17_out[7]) );
  INVX2TS U3311 ( .A(m17_out[7]), .Y(n2487) );
  INVX2TS U3312 ( .A(\alutwo/N324 ), .Y(n2457) );
  NOR3X2TS U3313 ( .A(alu2[1]), .B(alu2[0]), .C(n2457), .Y(n4710) );
  AOI22X1TS U3314 ( .A0(n3106), .A1(regeq_out[6]), .B0(n2452), .B1(
        regec_out[6]), .Y(n2440) );
  AOI22X1TS U3315 ( .A0(n3104), .A1(regep_out[6]), .B0(n2451), .B1(
        regea_out[6]), .Y(n2439) );
  NAND2X1TS U3316 ( .A(n2440), .B(n2439), .Y(m17_out[6]) );
  INVX2TS U3317 ( .A(m17_out[6]), .Y(n3504) );
  AOI22X1TS U3318 ( .A0(n3106), .A1(regeq_out[5]), .B0(n2452), .B1(
        regec_out[5]), .Y(n2442) );
  AOI22X1TS U3319 ( .A0(n3104), .A1(regep_out[5]), .B0(n2451), .B1(
        regea_out[5]), .Y(n2441) );
  NAND2X1TS U3320 ( .A(n2442), .B(n2441), .Y(m17_out[5]) );
  AOI22X1TS U3321 ( .A0(n3104), .A1(regep_out[4]), .B0(n2451), .B1(
        regea_out[4]), .Y(n2444) );
  AOI22X1TS U3322 ( .A0(n3106), .A1(regeq_out[4]), .B0(n2452), .B1(
        regec_out[4]), .Y(n2443) );
  NAND2X1TS U3323 ( .A(n2444), .B(n2443), .Y(m17_out[4]) );
  INVX2TS U3324 ( .A(m17_out[4]), .Y(n3456) );
  AOI22X1TS U3325 ( .A0(n3106), .A1(regeq_out[3]), .B0(n2452), .B1(
        regec_out[3]), .Y(n2446) );
  AOI22X1TS U3326 ( .A0(n3104), .A1(regep_out[3]), .B0(n2451), .B1(
        regea_out[3]), .Y(n2445) );
  NAND2X1TS U3327 ( .A(n2446), .B(n2445), .Y(m17_out[3]) );
  INVX2TS U3328 ( .A(m17_out[3]), .Y(n3446) );
  AOI22X1TS U3329 ( .A0(n3104), .A1(regep_out[2]), .B0(n2452), .B1(
        regec_out[2]), .Y(n2448) );
  AOI22X1TS U3330 ( .A0(n3106), .A1(regeq_out[2]), .B0(n2451), .B1(
        regea_out[2]), .Y(n2447) );
  NAND2X1TS U3331 ( .A(n2448), .B(n2447), .Y(m17_out[2]) );
  AOI22X1TS U3332 ( .A0(n3106), .A1(regeq_out[0]), .B0(n2452), .B1(
        regec_out[0]), .Y(n2450) );
  AOI22X1TS U3333 ( .A0(n3104), .A1(regep_out[0]), .B0(n2451), .B1(
        regea_out[0]), .Y(n2449) );
  NAND2X1TS U3334 ( .A(n2450), .B(n2449), .Y(m17_out[0]) );
  AOI22X1TS U3335 ( .A0(n3104), .A1(regep_out[1]), .B0(n2451), .B1(
        regea_out[1]), .Y(n2454) );
  AOI22X1TS U3336 ( .A0(n3106), .A1(regeq_out[1]), .B0(n2452), .B1(
        regec_out[1]), .Y(n2453) );
  NAND2X1TS U3337 ( .A(n2454), .B(n2453), .Y(m17_out[1]) );
  NAND2X1TS U3338 ( .A(n3504), .B(n3490), .Y(n2918) );
  NAND2X1TS U3339 ( .A(alu2[1]), .B(n2457), .Y(n4722) );
  INVX2TS U3340 ( .A(n4722), .Y(n3526) );
  AOI21X1TS U3341 ( .A0(n4710), .A1(n2918), .B0(n3526), .Y(n2486) );
  INVX2TS U3342 ( .A(n4710), .Y(n4660) );
  NAND2X1TS U3343 ( .A(m17_out[3]), .B(n2461), .Y(n2463) );
  NAND2X1TS U3344 ( .A(m17_out[5]), .B(n2465), .Y(n2468) );
  NAND2X1TS U3345 ( .A(m17_out[7]), .B(n2467), .Y(n2920) );
  OA21XLTS U3346 ( .A0(m17_out[7]), .A1(n2467), .B0(n2920), .Y(n2484) );
  INVX2TS U3347 ( .A(alu2[0]), .Y(n2922) );
  NAND2X1TS U3348 ( .A(\alutwo/N324 ), .B(alu2[1]), .Y(n2456) );
  NOR2X1TS U3349 ( .A(n2922), .B(n2456), .Y(n3493) );
  NAND2X1TS U3350 ( .A(n2457), .B(alu2[0]), .Y(n3503) );
  INVX2TS U3351 ( .A(n3507), .Y(m18_out[6]) );
  NOR2XLTS U3352 ( .A(regeb_out[5]), .B(n2458), .Y(n2474) );
  INVX2TS U3353 ( .A(n2474), .Y(m18_out[5]) );
  INVX2TS U3354 ( .A(n3459), .Y(m18_out[4]) );
  INVX2TS U3355 ( .A(n3339), .Y(m18_out[3]) );
  INVX2TS U3356 ( .A(n3311), .Y(m18_out[2]) );
  NOR2XLTS U3357 ( .A(regeb_out[1]), .B(n2458), .Y(n2471) );
  INVX2TS U3358 ( .A(n2471), .Y(m18_out[1]) );
  NAND2X1TS U3359 ( .A(n3303), .B(m17_out[1]), .Y(n2872) );
  AOI21X1TS U3360 ( .A0(m17_out[0]), .A1(m17_out[1]), .B0(n3309), .Y(n2878) );
  AOI21X1TS U3361 ( .A0(m18_out[1]), .A1(n2872), .B0(n2871), .Y(n2460) );
  INVX2TS U3362 ( .A(m17_out[2]), .Y(n3326) );
  NAND2X1TS U3363 ( .A(m17_out[0]), .B(m17_out[1]), .Y(n2459) );
  AOI21X1TS U3364 ( .A0(n3326), .A1(n2459), .B0(n2461), .Y(n3316) );
  NAND2X1TS U3365 ( .A(n2460), .B(n3316), .Y(n3318) );
  AOI21X1TS U3366 ( .A0(m18_out[2]), .A1(n3318), .B0(n3317), .Y(n2462) );
  OA21XLTS U3367 ( .A0(m17_out[3]), .A1(n2461), .B0(n2463), .Y(n3330) );
  NAND2X1TS U3368 ( .A(n2462), .B(n3330), .Y(n3332) );
  AOI21X1TS U3369 ( .A0(m18_out[3]), .A1(n3332), .B0(n3331), .Y(n2464) );
  AOI21X1TS U3370 ( .A0(n3456), .A1(n2463), .B0(n2465), .Y(n3448) );
  NAND2X1TS U3371 ( .A(n2464), .B(n3448), .Y(n3450) );
  AOI21X1TS U3372 ( .A0(m18_out[4]), .A1(n3450), .B0(n3449), .Y(n2466) );
  OA21XLTS U3373 ( .A0(m17_out[5]), .A1(n2465), .B0(n2468), .Y(n3385) );
  NAND2X1TS U3374 ( .A(n2466), .B(n3385), .Y(n3376) );
  AOI21X1TS U3375 ( .A0(m18_out[5]), .A1(n3376), .B0(n3375), .Y(n2469) );
  AOI21X1TS U3376 ( .A0(n3504), .A1(n2468), .B0(n2467), .Y(n3492) );
  NAND2X1TS U3377 ( .A(n2469), .B(n3492), .Y(n3495) );
  AOI21X1TS U3378 ( .A0(m18_out[6]), .A1(n3495), .B0(n3494), .Y(n2470) );
  NAND2X1TS U3379 ( .A(n2470), .B(n2484), .Y(n2921) );
  INVX2TS U3380 ( .A(n2456), .Y(n4696) );
  NAND2X1TS U3381 ( .A(n4696), .B(n2922), .Y(n3497) );
  OAI22X1TS U3382 ( .A0(n2487), .A1(n3503), .B0(n2479), .B1(n3497), .Y(n2478)
         );
  AOI21X1TS U3383 ( .A0(m18_out[0]), .A1(m17_out[0]), .B0(m17_out[1]), .Y(
        n2869) );
  AOI222XLTS U3384 ( .A0(m17_out[2]), .A1(m18_out[2]), .B0(m17_out[2]), .B1(
        n3320), .C0(m18_out[2]), .C1(n3320), .Y(n3333) );
  AOI222XLTS U3385 ( .A0(n3446), .A1(n3339), .B0(n3446), .B1(n3333), .C0(n3339), .C1(n3333), .Y(n2472) );
  NAND2X1TS U3386 ( .A(m17_out[4]), .B(n2472), .Y(n3451) );
  AOI21X1TS U3387 ( .A0(n3459), .A1(n3451), .B0(n3452), .Y(n2473) );
  NAND2X1TS U3388 ( .A(n2473), .B(m17_out[5]), .Y(n3373) );
  AOI21X1TS U3389 ( .A0(n2474), .A1(n3373), .B0(n3374), .Y(n3496) );
  AOI222XLTS U3390 ( .A0(n3496), .A1(m17_out[6]), .B0(n3496), .B1(m18_out[6]), 
        .C0(m17_out[6]), .C1(m18_out[6]), .Y(n2475) );
  NAND2X1TS U3391 ( .A(n2487), .B(n2475), .Y(n2937) );
  INVX2TS U3392 ( .A(n2937), .Y(n2477) );
  INVX2TS U3393 ( .A(alu2[1]), .Y(n2476) );
  INVX2TS U3394 ( .A(n4715), .Y(n4689) );
  OAI32X1TS U3395 ( .A0(n2478), .A1(n2936), .A2(n2477), .B0(n4689), .B1(n2478), 
        .Y(n2482) );
  NAND2X1TS U3396 ( .A(mux17[2]), .B(regeb_out[7]), .Y(n2480) );
  INVX2TS U3397 ( .A(n2480), .Y(m18_out[7]) );
  NAND2X1TS U3398 ( .A(alu2[0]), .B(n3526), .Y(n3501) );
  INVX2TS U3399 ( .A(n3497), .Y(n3499) );
  NOR2XLTS U3400 ( .A(n2936), .B(n4715), .Y(n3476) );
  AOI22X1TS U3401 ( .A0(n3499), .A1(n2479), .B0(n3476), .B1(n2937), .Y(n2481)
         );
  AOI32X1TS U3402 ( .A0(n2482), .A1(m18_out[7]), .A2(n3501), .B0(n2481), .B1(
        n2480), .Y(n2483) );
  AOI21X1TS U3403 ( .A0(n2484), .A1(n3493), .B0(n2483), .Y(n2485) );
  OAI221XLTS U3404 ( .A0(n2487), .A1(n2486), .B0(m17_out[7]), .B1(n3510), .C0(
        n2485), .Y(alutwo_out[7]) );
  AOI22X1TS U3405 ( .A0(n3125), .A1(srmt_out[12]), .B0(n3123), .B1(
        regms_out[12]), .Y(n2489) );
  AOI22X1TS U3406 ( .A0(n3124), .A1(reges0_out[12]), .B0(n2699), .B1(
        regres_out[12]), .Y(n2488) );
  NAND2X1TS U3407 ( .A(n2489), .B(n2488), .Y(n2519) );
  INVX2TS U3408 ( .A(n2519), .Y(n2525) );
  AOI22X1TS U3409 ( .A0(n3124), .A1(reges0_out[11]), .B0(n2699), .B1(
        regres_out[11]), .Y(n2490) );
  OAI2BB1X1TS U3410 ( .A0N(n3125), .A1N(srmt_out[11]), .B0(n2490), .Y(n2491)
         );
  AOI21X1TS U3411 ( .A0(n3123), .A1(regms_out[11]), .B0(n2491), .Y(n2902) );
  INVX2TS U3412 ( .A(n2902), .Y(n2907) );
  AOI22X1TS U3413 ( .A0(n3124), .A1(reges0_out[10]), .B0(n3123), .B1(
        regms_out[10]), .Y(n2493) );
  AOI22X1TS U3414 ( .A0(n3125), .A1(srmt_out[10]), .B0(n3122), .B1(
        regres_out[10]), .Y(n2492) );
  NAND2X1TS U3415 ( .A(n2493), .B(n2492), .Y(n2890) );
  INVX2TS U3416 ( .A(n2890), .Y(n2885) );
  NAND2X1TS U3417 ( .A(n2885), .B(n2883), .Y(n2735) );
  AOI21X1TS U3418 ( .A0(n2735), .A1(n3729), .B0(n3728), .Y(n2733) );
  INVX2TS U3419 ( .A(n2733), .Y(n2901) );
  AOI21X1TS U3420 ( .A0(n3729), .A1(n2907), .B0(n2901), .Y(n2520) );
  NAND2X1TS U3421 ( .A(n2525), .B(n2902), .Y(n2595) );
  INVX2TS U3422 ( .A(n2595), .Y(n2548) );
  NOR2X1TS U3423 ( .A(n2735), .B(n3357), .Y(n2948) );
  AOI21X1TS U3424 ( .A0(n2548), .A1(n2948), .B0(n2947), .Y(n2541) );
  AOI222X1TS U3425 ( .A0(ssrms0_out[12]), .A1(n2630), .B0(n2388), .B1(
        regms_out[12]), .C0(n3132), .C1(srmt_out[12]), .Y(n2531) );
  AOI222X1TS U3426 ( .A0(ssrms0_out[11]), .A1(n2630), .B0(n2388), .B1(
        regms_out[11]), .C0(n3132), .C1(srmt_out[11]), .Y(n2914) );
  AOI222X1TS U3427 ( .A0(ssrms0_out[10]), .A1(n2630), .B0(n2388), .B1(
        regms_out[10]), .C0(n3132), .C1(srmt_out[10]), .Y(n2897) );
  AOI21X1TS U3428 ( .A0(n2506), .A1(n2497), .B0(n2496), .Y(n2500) );
  NAND2X1TS U3429 ( .A(n2500), .B(n2900), .Y(n2888) );
  AOI21X1TS U3430 ( .A0(n2897), .A1(n2888), .B0(n2889), .Y(n2503) );
  NAND2X1TS U3431 ( .A(n2907), .B(n2502), .Y(n2526) );
  NAND2X1TS U3432 ( .A(n2503), .B(n2917), .Y(n2905) );
  AOI21X1TS U3433 ( .A0(n2914), .A1(n2905), .B0(n2906), .Y(n2504) );
  NAND2X1TS U3434 ( .A(n2504), .B(n2514), .Y(n2524) );
  AOI222XLTS U3435 ( .A0(n2507), .A1(n2506), .B0(n2507), .B1(n2505), .C0(n2506), .C1(n2505), .Y(n2508) );
  NAND2X1TS U3436 ( .A(n2508), .B(n2890), .Y(n2886) );
  AOI21X1TS U3437 ( .A0(n2897), .A1(n2886), .B0(n2887), .Y(n2509) );
  NAND2X1TS U3438 ( .A(n2509), .B(n2907), .Y(n2903) );
  AOI21X1TS U3439 ( .A0(n2914), .A1(n2903), .B0(n2904), .Y(n2510) );
  NAND2X1TS U3440 ( .A(n2510), .B(n2519), .Y(n2530) );
  NOR2BX1TS U3441 ( .AN(n2530), .B(n2529), .Y(n2512) );
  OAI22X1TS U3442 ( .A0(n2512), .A1(n3741), .B0(n3739), .B1(n2511), .Y(n2513)
         );
  OAI22X1TS U3443 ( .A0(n2531), .A1(n2515), .B0(n2514), .B1(n3748), .Y(n2516)
         );
  AOI21X1TS U3444 ( .A0(n2531), .A1(n2517), .B0(n2516), .Y(n2518) );
  OAI221XLTS U3445 ( .A0(n2525), .A1(n2520), .B0(n2519), .B1(n2541), .C0(n2518), .Y(aluone_out[12]) );
  AOI22X1TS U3446 ( .A0(n3123), .A1(regms_out[13]), .B0(n2699), .B1(
        regres_out[13]), .Y(n2521) );
  OAI2BB1X1TS U3447 ( .A0N(n3125), .A1N(srmt_out[13]), .B0(n2521), .Y(n2522)
         );
  AOI21X1TS U3448 ( .A0(n3124), .A1(reges0_out[13]), .B0(n2522), .Y(n2546) );
  AOI21X1TS U3449 ( .A0(n3729), .A1(n2595), .B0(n2901), .Y(n2542) );
  INVX2TS U3450 ( .A(n2546), .Y(n2545) );
  AOI222X1TS U3451 ( .A0(ssrms0_out[13]), .A1(n2630), .B0(n2388), .B1(
        regms_out[13]), .C0(n3132), .C1(srmt_out[13]), .Y(n2554) );
  AOI21X1TS U3452 ( .A0(n2531), .A1(n2524), .B0(n2523), .Y(n2528) );
  NAND2X1TS U3453 ( .A(n2545), .B(n2527), .Y(n2571) );
  NAND2X1TS U3454 ( .A(n2528), .B(n2536), .Y(n2550) );
  AOI21X1TS U3455 ( .A0(n2531), .A1(n2530), .B0(n2529), .Y(n2532) );
  NAND2X1TS U3456 ( .A(n2532), .B(n2545), .Y(n2553) );
  NOR2BX1TS U3457 ( .AN(n2553), .B(n2552), .Y(n2534) );
  OAI22X1TS U3458 ( .A0(n2534), .A1(n3741), .B0(n3739), .B1(n2533), .Y(n2535)
         );
  OAI22X1TS U3459 ( .A0(n2554), .A1(n2537), .B0(n2536), .B1(n3748), .Y(n2538)
         );
  AOI21X1TS U3460 ( .A0(n2554), .A1(n2539), .B0(n2538), .Y(n2540) );
  OAI221XLTS U3461 ( .A0(n2546), .A1(n2542), .B0(n2545), .B1(n2541), .C0(n2540), .Y(aluone_out[13]) );
  AOI22X1TS U3462 ( .A0(n3123), .A1(regms_out[14]), .B0(n3122), .B1(
        regres_out[14]), .Y(n2544) );
  AOI22X1TS U3463 ( .A0(n3124), .A1(reges0_out[14]), .B0(n3125), .B1(
        srmt_out[14]), .Y(n2543) );
  NAND2X1TS U3464 ( .A(n2544), .B(n2543), .Y(n2564) );
  INVX2TS U3465 ( .A(n2564), .Y(n2570) );
  OAI32X1TS U3466 ( .A0(n2901), .A1(n2595), .A2(n2545), .B0(n3729), .B1(n2901), 
        .Y(n2565) );
  NAND2X1TS U3467 ( .A(n2570), .B(n2546), .Y(n2596) );
  INVX2TS U3468 ( .A(n2596), .Y(n2547) );
  AOI222X1TS U3469 ( .A0(ssrms0_out[14]), .A1(n2630), .B0(n2388), .B1(
        regms_out[14]), .C0(n3132), .C1(srmt_out[14]), .Y(n2576) );
  AOI21X1TS U3470 ( .A0(n2554), .A1(n2550), .B0(n2549), .Y(n2551) );
  NAND2X1TS U3471 ( .A(n2551), .B(n2559), .Y(n2569) );
  AOI21X1TS U3472 ( .A0(n2554), .A1(n2553), .B0(n2552), .Y(n2555) );
  NAND2X1TS U3473 ( .A(n2555), .B(n2564), .Y(n2575) );
  NOR2BX1TS U3474 ( .AN(n2575), .B(n2574), .Y(n2557) );
  OAI22X1TS U3475 ( .A0(n2557), .A1(n3741), .B0(n3739), .B1(n2556), .Y(n2558)
         );
  OAI22X1TS U3476 ( .A0(n2576), .A1(n2560), .B0(n2559), .B1(n3748), .Y(n2561)
         );
  AOI21X1TS U3477 ( .A0(n2576), .A1(n2562), .B0(n2561), .Y(n2563) );
  OAI221XLTS U3478 ( .A0(n2570), .A1(n2565), .B0(n2564), .B1(n2586), .C0(n2563), .Y(aluone_out[14]) );
  AOI22X1TS U3479 ( .A0(n3124), .A1(reges0_out[15]), .B0(n3123), .B1(
        regms_out[15]), .Y(n2566) );
  OAI2BB1X1TS U3480 ( .A0N(n3125), .A1N(srmt_out[15]), .B0(n2566), .Y(n2567)
         );
  AOI21X1TS U3481 ( .A0(n3122), .A1(regres_out[15]), .B0(n2567), .Y(n2966) );
  OAI32X1TS U3482 ( .A0(n2901), .A1(n2595), .A2(n2596), .B0(n3729), .B1(n2901), 
        .Y(n2965) );
  INVX2TS U3483 ( .A(n2966), .Y(n2597) );
  AOI222X1TS U3484 ( .A0(ssrms0_out[15]), .A1(n2630), .B0(n2388), .B1(
        regms_out[15]), .C0(n3132), .C1(srmt_out[15]), .Y(n2610) );
  AOI21X1TS U3485 ( .A0(n2576), .A1(n2569), .B0(n2568), .Y(n2573) );
  NAND2X1TS U3486 ( .A(n2597), .B(n2572), .Y(n2601) );
  NAND2X1TS U3487 ( .A(n2573), .B(n2581), .Y(n2599) );
  AOI21X1TS U3488 ( .A0(n2576), .A1(n2575), .B0(n2574), .Y(n2577) );
  NAND2X1TS U3489 ( .A(n2577), .B(n2597), .Y(n2609) );
  NOR2BX1TS U3490 ( .AN(n2609), .B(n2608), .Y(n2579) );
  OAI22X1TS U3491 ( .A0(n2579), .A1(n3741), .B0(n3739), .B1(n2578), .Y(n2580)
         );
  OAI22X1TS U3492 ( .A0(n2610), .A1(n2582), .B0(n2581), .B1(n3748), .Y(n2583)
         );
  AOI21X1TS U3493 ( .A0(n2610), .A1(n2584), .B0(n2583), .Y(n2585) );
  OAI221XLTS U3494 ( .A0(n2966), .A1(n2965), .B0(n2597), .B1(n2586), .C0(n2585), .Y(aluone_out[15]) );
  AOI22X1TS U3495 ( .A0(n3124), .A1(reges0_out[19]), .B0(n3123), .B1(
        regms_out[19]), .Y(n2587) );
  OAI2BB1X1TS U3496 ( .A0N(n3125), .A1N(srmt_out[19]), .B0(n2587), .Y(n2588)
         );
  AOI21X1TS U3497 ( .A0(n3122), .A1(regres_out[19]), .B0(n2588), .Y(n3005) );
  AOI22X1TS U3498 ( .A0(n3125), .A1(srmt_out[18]), .B0(n3123), .B1(
        regms_out[18]), .Y(n2590) );
  AOI22X1TS U3499 ( .A0(n3124), .A1(reges0_out[18]), .B0(n2699), .B1(
        regres_out[18]), .Y(n2589) );
  NAND2X1TS U3500 ( .A(n2590), .B(n2589), .Y(n3001) );
  AOI22X1TS U3501 ( .A0(n3124), .A1(reges0_out[17]), .B0(n3123), .B1(
        regms_out[17]), .Y(n2591) );
  OAI2BB1X1TS U3502 ( .A0N(n3125), .A1N(srmt_out[17]), .B0(n2591), .Y(n2592)
         );
  AOI21X1TS U3503 ( .A0(n3122), .A1(regres_out[17]), .B0(n2592), .Y(n2950) );
  INVX2TS U3504 ( .A(n2950), .Y(n2998) );
  AOI22X1TS U3505 ( .A0(n3124), .A1(reges0_out[16]), .B0(n3122), .B1(
        regres_out[16]), .Y(n2594) );
  AOI22X1TS U3506 ( .A0(n3125), .A1(srmt_out[16]), .B0(n3123), .B1(
        regms_out[16]), .Y(n2593) );
  NAND2X1TS U3507 ( .A(n2594), .B(n2593), .Y(n2974) );
  INVX2TS U3508 ( .A(n3005), .Y(n2629) );
  AOI222X1TS U3509 ( .A0(ssrms0_out[19]), .A1(n2630), .B0(n2388), .B1(
        regms_out[19]), .C0(n3132), .C1(srmt_out[19]), .Y(n2640) );
  AOI222X1TS U3510 ( .A0(ssrms0_out[18]), .A1(n2630), .B0(n2388), .B1(
        regms_out[18]), .C0(n3132), .C1(srmt_out[18]), .Y(n2996) );
  AOI222X1TS U3511 ( .A0(ssrms0_out[17]), .A1(n2630), .B0(n2388), .B1(
        regms_out[17]), .C0(n3132), .C1(srmt_out[17]), .Y(n2961) );
  AOI222XLTS U3512 ( .A0(ssrms0_out[16]), .A1(n2630), .B0(n2388), .B1(
        regms_out[16]), .C0(n3132), .C1(srmt_out[16]), .Y(n2981) );
  AOI21X1TS U3513 ( .A0(n2610), .A1(n2599), .B0(n2598), .Y(n2600) );
  NAND2X1TS U3514 ( .A(n2600), .B(n2984), .Y(n2972) );
  AOI21X1TS U3515 ( .A0(n2981), .A1(n2972), .B0(n2973), .Y(n2603) );
  INVX2TS U3516 ( .A(n2974), .Y(n2969) );
  NAND2X1TS U3517 ( .A(n2998), .B(n2602), .Y(n2605) );
  NAND2X1TS U3518 ( .A(n2603), .B(n2964), .Y(n2953) );
  AOI21X1TS U3519 ( .A0(n2961), .A1(n2953), .B0(n2954), .Y(n2604) );
  NAND2X1TS U3520 ( .A(n2604), .B(n2992), .Y(n2985) );
  AOI21X1TS U3521 ( .A0(n2996), .A1(n2985), .B0(n2986), .Y(n2607) );
  NOR2BX1TS U3522 ( .AN(n3001), .B(n2605), .Y(n2606) );
  NAND2X1TS U3523 ( .A(n2629), .B(n2606), .Y(n2634) );
  NAND2X1TS U3524 ( .A(n2607), .B(n2618), .Y(n2632) );
  AOI21X1TS U3525 ( .A0(n2610), .A1(n2609), .B0(n2608), .Y(n2611) );
  NAND2X1TS U3526 ( .A(n2611), .B(n2974), .Y(n2970) );
  OAI21XLTS U3527 ( .A0(n2981), .A1(n2971), .B0(n2970), .Y(n2612) );
  NAND2X1TS U3528 ( .A(n2998), .B(n2612), .Y(n2951) );
  AOI21X1TS U3529 ( .A0(n2961), .A1(n2951), .B0(n2952), .Y(n2613) );
  NAND2X1TS U3530 ( .A(n2613), .B(n3001), .Y(n2988) );
  AOI21X1TS U3531 ( .A0(n2996), .A1(n2988), .B0(n2987), .Y(n2614) );
  NAND2X1TS U3532 ( .A(n2614), .B(n2629), .Y(n2639) );
  NOR2BX1TS U3533 ( .AN(n2639), .B(n2638), .Y(n2616) );
  OAI22X1TS U3534 ( .A0(n2616), .A1(n3741), .B0(n3739), .B1(n2615), .Y(n2617)
         );
  OAI22X1TS U3535 ( .A0(n2640), .A1(n2619), .B0(n2618), .B1(n3748), .Y(n2620)
         );
  AOI21X1TS U3536 ( .A0(n2640), .A1(n2621), .B0(n2620), .Y(n2622) );
  OAI221XLTS U3537 ( .A0(n3005), .A1(n3004), .B0(n2629), .B1(n3002), .C0(n2622), .Y(aluone_out[19]) );
  AOI22X1TS U3538 ( .A0(n3124), .A1(reges0_out[22]), .B0(n3123), .B1(
        regms_out[22]), .Y(n2624) );
  AOI22X1TS U3539 ( .A0(n3125), .A1(srmt_out[22]), .B0(n3122), .B1(
        regres_out[22]), .Y(n2623) );
  NAND2X1TS U3540 ( .A(n2624), .B(n2623), .Y(n2652) );
  INVX2TS U3541 ( .A(n2652), .Y(n2658) );
  AOI22X1TS U3542 ( .A0(n3124), .A1(reges0_out[21]), .B0(n2699), .B1(
        regres_out[21]), .Y(n2625) );
  OAI2BB1X1TS U3543 ( .A0N(n3125), .A1N(srmt_out[21]), .B0(n2625), .Y(n2626)
         );
  AOI21X1TS U3544 ( .A0(n3123), .A1(regms_out[21]), .B0(n2626), .Y(n3025) );
  INVX2TS U3545 ( .A(n3025), .Y(n3030) );
  AOI22X1TS U3546 ( .A0(n3125), .A1(srmt_out[20]), .B0(n3122), .B1(
        regres_out[20]), .Y(n2628) );
  AOI22X1TS U3547 ( .A0(n3124), .A1(reges0_out[20]), .B0(n3123), .B1(
        regms_out[20]), .Y(n2627) );
  NAND2X1TS U3548 ( .A(n2628), .B(n2627), .Y(n3012) );
  AOI21X1TS U3549 ( .A0(n3729), .A1(n3030), .B0(n3023), .Y(n2653) );
  NAND2X1TS U3550 ( .A(n2658), .B(n3025), .Y(n2678) );
  AOI222X1TS U3551 ( .A0(ssrms0_out[22]), .A1(n2630), .B0(n2388), .B1(
        regms_out[22]), .C0(n3132), .C1(srmt_out[22]), .Y(n2663) );
  AOI222XLTS U3552 ( .A0(ssrms0_out[21]), .A1(n2630), .B0(n2388), .B1(
        regms_out[21]), .C0(n3132), .C1(srmt_out[21]), .Y(n3037) );
  AOI222XLTS U3553 ( .A0(ssrms0_out[20]), .A1(n2630), .B0(n2388), .B1(
        regms_out[20]), .C0(n3132), .C1(srmt_out[20]), .Y(n3019) );
  AOI21X1TS U3554 ( .A0(n2640), .A1(n2632), .B0(n2631), .Y(n2633) );
  NAND2X1TS U3555 ( .A(n2633), .B(n3022), .Y(n3010) );
  AOI21X1TS U3556 ( .A0(n3019), .A1(n3010), .B0(n3011), .Y(n2636) );
  INVX2TS U3557 ( .A(n3012), .Y(n3007) );
  NAND2X1TS U3558 ( .A(n3030), .B(n2635), .Y(n2659) );
  NAND2X1TS U3559 ( .A(n2636), .B(n3040), .Y(n3028) );
  AOI21X1TS U3560 ( .A0(n3037), .A1(n3028), .B0(n3029), .Y(n2637) );
  NAND2X1TS U3561 ( .A(n2637), .B(n2647), .Y(n2657) );
  AOI21X1TS U3562 ( .A0(n2640), .A1(n2639), .B0(n2638), .Y(n2641) );
  NAND2X1TS U3563 ( .A(n2641), .B(n3012), .Y(n3008) );
  OAI21XLTS U3564 ( .A0(n3019), .A1(n3009), .B0(n3008), .Y(n2642) );
  NAND2X1TS U3565 ( .A(n3030), .B(n2642), .Y(n3026) );
  OAI21XLTS U3566 ( .A0(n3037), .A1(n3027), .B0(n3026), .Y(n2643) );
  NAND2X1TS U3567 ( .A(n2652), .B(n2643), .Y(n2661) );
  NOR2BX1TS U3568 ( .AN(n2661), .B(n2662), .Y(n2645) );
  OAI22X1TS U3569 ( .A0(n2645), .A1(n3741), .B0(n3739), .B1(n2644), .Y(n2646)
         );
  OAI22X1TS U3570 ( .A0(n2663), .A1(n2648), .B0(n2647), .B1(n3748), .Y(n2649)
         );
  AOI21X1TS U3571 ( .A0(n2663), .A1(n2650), .B0(n2649), .Y(n2651) );
  OAI221XLTS U3572 ( .A0(n2658), .A1(n2653), .B0(n2652), .B1(n2673), .C0(n2651), .Y(aluone_out[22]) );
  AOI22X1TS U3573 ( .A0(n3124), .A1(reges0_out[23]), .B0(n3122), .B1(
        regres_out[23]), .Y(n2654) );
  OAI2BB1X1TS U3574 ( .A0N(n3125), .A1N(srmt_out[23]), .B0(n2654), .Y(n2655)
         );
  AOI21X1TS U3575 ( .A0(n2702), .A1(regms_out[23]), .B0(n2655), .Y(n2675) );
  AOI21X1TS U3576 ( .A0(n3729), .A1(n2678), .B0(n3023), .Y(n2674) );
  INVX2TS U3577 ( .A(n2675), .Y(n2682) );
  AOI222X1TS U3578 ( .A0(ssrms0_out[23]), .A1(n2630), .B0(n2388), .B1(
        regms_out[23]), .C0(n3132), .C1(srmt_out[23]), .Y(n2687) );
  AOI21X1TS U3579 ( .A0(n2663), .A1(n2657), .B0(n2656), .Y(n2660) );
  NAND2X1TS U3580 ( .A(n2660), .B(n2668), .Y(n2681) );
  OAI21XLTS U3581 ( .A0(n2663), .A1(n2662), .B0(n2661), .Y(n2664) );
  NAND2X1TS U3582 ( .A(n2682), .B(n2664), .Y(n2686) );
  NOR2BX1TS U3583 ( .AN(n2686), .B(n2685), .Y(n2666) );
  OAI22X1TS U3584 ( .A0(n2666), .A1(n3741), .B0(n3739), .B1(n2665), .Y(n2667)
         );
  OAI22X1TS U3585 ( .A0(n2687), .A1(n2669), .B0(n2668), .B1(n3748), .Y(n2670)
         );
  AOI21X1TS U3586 ( .A0(n2687), .A1(n2671), .B0(n2670), .Y(n2672) );
  OAI221XLTS U3587 ( .A0(n2675), .A1(n2674), .B0(n2682), .B1(n2673), .C0(n2672), .Y(aluone_out[23]) );
  AOI22X1TS U3588 ( .A0(n3124), .A1(reges0_out[24]), .B0(n3125), .B1(
        srmt_out[24]), .Y(n2677) );
  AOI22X1TS U3589 ( .A0(n3123), .A1(regms_out[24]), .B0(n3122), .B1(
        regres_out[24]), .Y(n2676) );
  NAND2X1TS U3590 ( .A(n2677), .B(n2676), .Y(n2697) );
  INVX2TS U3591 ( .A(n2697), .Y(n2705) );
  NAND2X1TS U3592 ( .A(n2705), .B(n2679), .Y(n2732) );
  AOI222X1TS U3593 ( .A0(n2388), .A1(regms_out[24]), .B0(n2630), .B1(
        ssrms0_out[24]), .C0(n3132), .C1(srmt_out[24]), .Y(n2711) );
  AOI21X1TS U3594 ( .A0(n2687), .A1(n2681), .B0(n2680), .Y(n2684) );
  NAND2X1TS U3595 ( .A(n2684), .B(n2692), .Y(n2704) );
  AOI21X1TS U3596 ( .A0(n2687), .A1(n2686), .B0(n2685), .Y(n2688) );
  NAND2X1TS U3597 ( .A(n2688), .B(n2697), .Y(n2710) );
  NOR2BX1TS U3598 ( .AN(n2710), .B(n2709), .Y(n2690) );
  OAI22X1TS U3599 ( .A0(n2690), .A1(n3741), .B0(n3739), .B1(n2689), .Y(n2691)
         );
  OAI22X1TS U3600 ( .A0(n2711), .A1(n2693), .B0(n2692), .B1(n3748), .Y(n2694)
         );
  AOI21X1TS U3601 ( .A0(n2711), .A1(n2695), .B0(n2694), .Y(n2696) );
  OAI221XLTS U3602 ( .A0(n2705), .A1(n2698), .B0(n2697), .B1(n2721), .C0(n2696), .Y(aluone_out[24]) );
  AOI22X1TS U3603 ( .A0(n3124), .A1(reges0_out[25]), .B0(n2699), .B1(
        regres_out[25]), .Y(n2700) );
  OAI2BB1X1TS U3604 ( .A0N(n3125), .A1N(srmt_out[25]), .B0(n2700), .Y(n2701)
         );
  AOI21X1TS U3605 ( .A0(n2702), .A1(regms_out[25]), .B0(n2701), .Y(n3044) );
  AOI21X1TS U3606 ( .A0(n3729), .A1(n2732), .B0(n3023), .Y(n3043) );
  INVX2TS U3607 ( .A(n3044), .Y(n2728) );
  AOI222X1TS U3608 ( .A0(n2388), .A1(regms_out[25]), .B0(n2630), .B1(
        ssrms0_out[25]), .C0(n3132), .C1(srmt_out[25]), .Y(n2746) );
  AOI21X1TS U3609 ( .A0(n2711), .A1(n2704), .B0(n2703), .Y(n2708) );
  NAND2X1TS U3610 ( .A(n2728), .B(n2707), .Y(n2740) );
  NAND2X1TS U3611 ( .A(n2708), .B(n2716), .Y(n2738) );
  AOI21X1TS U3612 ( .A0(n2711), .A1(n2710), .B0(n2709), .Y(n2712) );
  NAND2X1TS U3613 ( .A(n2712), .B(n2728), .Y(n2744) );
  NOR2BX1TS U3614 ( .AN(n2744), .B(n2745), .Y(n2714) );
  OAI22X1TS U3615 ( .A0(n2714), .A1(n3741), .B0(n3739), .B1(n2713), .Y(n2715)
         );
  OAI22X1TS U3616 ( .A0(n2746), .A1(n2717), .B0(n2716), .B1(n3748), .Y(n2718)
         );
  AOI21X1TS U3617 ( .A0(n2746), .A1(n2719), .B0(n2718), .Y(n2720) );
  OAI221XLTS U3618 ( .A0(n3044), .A1(n3043), .B0(n2728), .B1(n2721), .C0(n2720), .Y(aluone_out[25]) );
  AOI22X1TS U3619 ( .A0(n3124), .A1(reges0_out[28]), .B0(n3125), .B1(
        srmt_out[28]), .Y(n2723) );
  AOI22X1TS U3620 ( .A0(n3123), .A1(regms_out[28]), .B0(n3122), .B1(
        regres_out[28]), .Y(n2722) );
  NAND2X1TS U3621 ( .A(n2723), .B(n2722), .Y(n2758) );
  INVX2TS U3622 ( .A(n2758), .Y(n2765) );
  AOI22X1TS U3623 ( .A0(n3123), .A1(regms_out[27]), .B0(n3122), .B1(
        regres_out[27]), .Y(n2724) );
  OAI2BB1X1TS U3624 ( .A0N(n3125), .A1N(srmt_out[27]), .B0(n2724), .Y(n2725)
         );
  AOI21X1TS U3625 ( .A0(n3124), .A1(reges0_out[27]), .B0(n2725), .Y(n3064) );
  INVX2TS U3626 ( .A(n3064), .Y(n3069) );
  AOI22X1TS U3627 ( .A0(n3125), .A1(srmt_out[26]), .B0(n3122), .B1(
        regres_out[26]), .Y(n2727) );
  AOI22X1TS U3628 ( .A0(n3124), .A1(reges0_out[26]), .B0(n3123), .B1(
        regms_out[26]), .Y(n2726) );
  NAND2X1TS U3629 ( .A(n2727), .B(n2726), .Y(n3051) );
  AOI21X1TS U3630 ( .A0(n3729), .A1(n3069), .B0(n3062), .Y(n2759) );
  AOI222X1TS U3631 ( .A0(n2388), .A1(regms_out[28]), .B0(n2630), .B1(
        ssrms0_out[28]), .C0(n3132), .C1(srmt_out[28]), .Y(n2771) );
  AOI222XLTS U3632 ( .A0(n2388), .A1(regms_out[27]), .B0(n2630), .B1(
        ssrms0_out[27]), .C0(n3132), .C1(srmt_out[27]), .Y(n3076) );
  AOI222XLTS U3633 ( .A0(n2388), .A1(regms_out[26]), .B0(n2630), .B1(
        ssrms0_out[26]), .C0(n3132), .C1(srmt_out[26]), .Y(n3058) );
  AOI21X1TS U3634 ( .A0(n2746), .A1(n2738), .B0(n2737), .Y(n2739) );
  NAND2X1TS U3635 ( .A(n2739), .B(n3061), .Y(n3049) );
  AOI21X1TS U3636 ( .A0(n3058), .A1(n3049), .B0(n3050), .Y(n2742) );
  INVX2TS U3637 ( .A(n3051), .Y(n3046) );
  NAND2X1TS U3638 ( .A(n3069), .B(n2741), .Y(n2766) );
  NAND2X1TS U3639 ( .A(n2742), .B(n3079), .Y(n3067) );
  AOI21X1TS U3640 ( .A0(n3076), .A1(n3067), .B0(n3068), .Y(n2743) );
  NAND2X1TS U3641 ( .A(n2743), .B(n2753), .Y(n2764) );
  OAI21XLTS U3642 ( .A0(n2746), .A1(n2745), .B0(n2744), .Y(n2747) );
  NAND2X1TS U3643 ( .A(n3051), .B(n2747), .Y(n3047) );
  OAI21XLTS U3644 ( .A0(n3058), .A1(n3048), .B0(n3047), .Y(n2748) );
  NAND2X1TS U3645 ( .A(n3069), .B(n2748), .Y(n3065) );
  OAI21XLTS U3646 ( .A0(n3076), .A1(n3066), .B0(n3065), .Y(n2749) );
  NAND2X1TS U3647 ( .A(n2758), .B(n2749), .Y(n2770) );
  NOR2BX1TS U3648 ( .AN(n2770), .B(n2769), .Y(n2751) );
  OAI22X1TS U3649 ( .A0(n2751), .A1(n3741), .B0(n3739), .B1(n2750), .Y(n2752)
         );
  OAI22X1TS U3650 ( .A0(n2771), .A1(n2754), .B0(n2753), .B1(n3748), .Y(n2755)
         );
  AOI21X1TS U3651 ( .A0(n2771), .A1(n2756), .B0(n2755), .Y(n2757) );
  OAI221XLTS U3652 ( .A0(n2765), .A1(n2759), .B0(n2758), .B1(n2781), .C0(n2757), .Y(aluone_out[28]) );
  AOI22X1TS U3653 ( .A0(n3124), .A1(reges0_out[29]), .B0(n3123), .B1(
        regms_out[29]), .Y(n2760) );
  OAI2BB1X1TS U3654 ( .A0N(n3125), .A1N(srmt_out[29]), .B0(n2760), .Y(n2761)
         );
  AOI21X1TS U3655 ( .A0(n3122), .A1(regres_out[29]), .B0(n2761), .Y(n3085) );
  AOI21X1TS U3656 ( .A0(n3729), .A1(n2762), .B0(n2901), .Y(n3084) );
  INVX2TS U3657 ( .A(n3085), .Y(n2782) );
  AOI222X1TS U3658 ( .A0(n2388), .A1(regms_out[29]), .B0(n2630), .B1(
        ssrms0_out[29]), .C0(n3132), .C1(srmt_out[29]), .Y(n3092) );
  AOI21X1TS U3659 ( .A0(n2771), .A1(n2764), .B0(n2763), .Y(n2768) );
  NAND2X1TS U3660 ( .A(n2782), .B(n2767), .Y(n3129) );
  NAND2X1TS U3661 ( .A(n2768), .B(n2776), .Y(n3091) );
  AOI21X1TS U3662 ( .A0(n2771), .A1(n2770), .B0(n2769), .Y(n2772) );
  NAND2X1TS U3663 ( .A(n2772), .B(n2782), .Y(n3087) );
  NOR2BX1TS U3664 ( .AN(n3087), .B(n3088), .Y(n2774) );
  OAI22X1TS U3665 ( .A0(n2774), .A1(n3741), .B0(n3739), .B1(n2773), .Y(n2775)
         );
  OAI22X1TS U3666 ( .A0(n3092), .A1(n2777), .B0(n2776), .B1(n3748), .Y(n2778)
         );
  AOI21X1TS U3667 ( .A0(n3092), .A1(n2779), .B0(n2778), .Y(n2780) );
  OAI221XLTS U3668 ( .A0(n3085), .A1(n3084), .B0(n2782), .B1(n2781), .C0(n2780), .Y(aluone_out[29]) );
  INVX2TS U3669 ( .A(mux19), .Y(n4610) );
  INVX2TS U3670 ( .A(n4610), .Y(n4612) );
  AO22X1TS U3671 ( .A0(n4612), .A1(regmc_out[0]), .B0(n4610), .B1(regma_out[0]), .Y(m19_out[0]) );
  AO22XLTS U3672 ( .A0(n4612), .A1(regmc_out[12]), .B0(n4610), .B1(
        regma_out[12]), .Y(m19_out[12]) );
  AO22XLTS U3673 ( .A0(n4612), .A1(regmc_out[15]), .B0(n4610), .B1(
        regma_out[15]), .Y(m19_out[15]) );
  AO22XLTS U3674 ( .A0(n4612), .A1(regmc_out[16]), .B0(n4610), .B1(
        regma_out[16]), .Y(m19_out[16]) );
  AO22XLTS U3675 ( .A0(n4612), .A1(regmc_out[17]), .B0(n4610), .B1(
        regma_out[17]), .Y(m19_out[17]) );
  AO22XLTS U3676 ( .A0(n4612), .A1(regmc_out[18]), .B0(n4610), .B1(
        regma_out[18]), .Y(m19_out[18]) );
  AO22XLTS U3677 ( .A0(n4612), .A1(regmc_out[19]), .B0(n4610), .B1(
        regma_out[19]), .Y(m19_out[19]) );
  AO22XLTS U3678 ( .A0(n4612), .A1(regmc_out[20]), .B0(n4610), .B1(
        regma_out[20]), .Y(m19_out[20]) );
  AO22XLTS U3679 ( .A0(n4612), .A1(regmc_out[21]), .B0(n4610), .B1(
        regma_out[21]), .Y(m19_out[21]) );
  AO22X1TS U3680 ( .A0(n4612), .A1(regmc_out[22]), .B0(n4610), .B1(
        regma_out[22]), .Y(m19_out[22]) );
  INVX2TS U3681 ( .A(mux15), .Y(n2783) );
  AO22XLTS U3682 ( .A0(mux15), .A1(regindex_out[5]), .B0(n2783), .B1(rf_rab[5]), .Y(m15_out[5]) );
  NOR2XLTS U3683 ( .A(n4784), .B(n2783), .Y(m15_out[4]) );
  NOR2XLTS U3684 ( .A(n4773), .B(n2783), .Y(m15_out[3]) );
  NOR2BX1TS U3685 ( .AN(regindex_out[2]), .B(n2783), .Y(m15_out[2]) );
  AO22XLTS U3686 ( .A0(mux15), .A1(regindex_out[1]), .B0(n2783), .B1(rf_rab[1]), .Y(m15_out[1]) );
  AO22XLTS U3687 ( .A0(mux15), .A1(regindex_out[0]), .B0(n2783), .B1(rf_rab[0]), .Y(m15_out[0]) );
  INVX2TS U3688 ( .A(ssrms0_out[16]), .Y(n4166) );
  INVX2TS U3689 ( .A(ssrms0_out[17]), .Y(n4147) );
  INVX2TS U3690 ( .A(ssrms0_out[18]), .Y(n4137) );
  INVX2TS U3691 ( .A(ssrms0_out[19]), .Y(n4127) );
  NAND4XLTS U3692 ( .A(n4166), .B(n4147), .C(n4137), .D(n4127), .Y(n3794) );
  NOR4XLTS U3693 ( .A(ssrms0_out[20]), .B(ssrms0_out[21]), .C(ssrms0_out[22]), 
        .D(n3794), .Y(n3811) );
  INVX2TS U3694 ( .A(ssrms0_out[12]), .Y(n4196) );
  INVX2TS U3695 ( .A(ssrms0_out[13]), .Y(n4189) );
  INVX2TS U3696 ( .A(ssrms0_out[14]), .Y(n4182) );
  INVX2TS U3697 ( .A(ssrms0_out[15]), .Y(n4175) );
  NAND4XLTS U3698 ( .A(n4196), .B(n4189), .C(n4182), .D(n4175), .Y(n3790) );
  NOR2XLTS U3699 ( .A(ssrms0_out[11]), .B(n3790), .Y(n3810) );
  NAND2X1TS U3700 ( .A(n3811), .B(n3810), .Y(n2798) );
  NOR2XLTS U3701 ( .A(ssrms0_out[10]), .B(n2798), .Y(n2793) );
  INVX2TS U3702 ( .A(ssrms0_out[9]), .Y(n4220) );
  NOR3XLTS U3703 ( .A(ssrms0_out[8]), .B(ssrms0_out[9]), .C(ssrms0_out[10]), 
        .Y(n3812) );
  NOR2XLTS U3704 ( .A(ssrms0_out[6]), .B(ssrms0_out[7]), .Y(n2792) );
  NAND4BXLTS U3705 ( .AN(n2798), .B(n3812), .C(n2792), .D(n4257), .Y(n2785) );
  INVX2TS U3706 ( .A(ssrms0_out[3]), .Y(n4276) );
  NAND2X1TS U3707 ( .A(n4286), .B(n4276), .Y(n2786) );
  INVX2TS U3708 ( .A(ssrms0_out[4]), .Y(n4266) );
  OAI32X1TS U3709 ( .A0(n2785), .A1(ssrms0_out[1]), .A2(n2786), .B0(n4266), 
        .B1(n2785), .Y(n2784) );
  AOI31XLTS U3710 ( .A0(ssrms0_out[8]), .A1(n2793), .A2(n4220), .B0(n2784), 
        .Y(n2804) );
  NOR2XLTS U3711 ( .A(ssrms0_out[4]), .B(n2785), .Y(n3793) );
  INVX2TS U3712 ( .A(n2786), .Y(n2791) );
  INVX2TS U3713 ( .A(ssrms0_out[20]), .Y(n4106) );
  INVX2TS U3714 ( .A(ssrms0_out[21]), .Y(n4100) );
  OAI211XLTS U3715 ( .A0(ssrms0_out[16]), .A1(ssrms0_out[17]), .B0(n4127), 
        .C0(n4137), .Y(n2787) );
  AOI31XLTS U3716 ( .A0(n4106), .A1(n4100), .A2(n2787), .B0(ssrms0_out[22]), 
        .Y(n2790) );
  INVX2TS U3717 ( .A(n3811), .Y(n3789) );
  NAND2X1TS U3718 ( .A(n4182), .B(n4175), .Y(n2788) );
  AOI211XLTS U3719 ( .A0(n4196), .A1(n4189), .B0(n3789), .C0(n2788), .Y(n2789)
         );
  AOI211XLTS U3720 ( .A0(n3793), .A1(n2791), .B0(n2790), .C0(n2789), .Y(n2795)
         );
  AOI32X1TS U3721 ( .A0(ssrms0_out[5]), .A1(n2793), .A2(n2792), .B0(
        ssrms0_out[9]), .B1(n2793), .Y(n2794) );
  AOI31XLTS U3722 ( .A0(n2804), .A1(n2795), .A2(n2794), .B0(ssrms0_out[23]), 
        .Y(pe_out[1]) );
  OAI21XLTS U3723 ( .A0(ssrms0_out[13]), .A1(n4196), .B0(n4182), .Y(n2796) );
  AOI31XLTS U3724 ( .A0(n3811), .A1(n4175), .A2(n2796), .B0(ssrms0_out[22]), 
        .Y(n2803) );
  OAI21XLTS U3725 ( .A0(ssrms0_out[17]), .A1(n4166), .B0(n4137), .Y(n2797) );
  AOI21X1TS U3726 ( .A0(n4127), .A1(n2797), .B0(ssrms0_out[20]), .Y(n2800) );
  INVX2TS U3727 ( .A(ssrms0_out[7]), .Y(n4239) );
  AOI31XLTS U3728 ( .A0(ssrms0_out[6]), .A1(n4220), .A2(n4239), .B0(
        ssrms0_out[10]), .Y(n2799) );
  OAI22X1TS U3729 ( .A0(ssrms0_out[21]), .A1(n2800), .B0(n2799), .B1(n2798), 
        .Y(n2801) );
  AOI31XLTS U3730 ( .A0(ssrms0_out[2]), .A1(n3793), .A2(n4276), .B0(n2801), 
        .Y(n2802) );
  AOI31XLTS U3731 ( .A0(n2804), .A1(n2803), .A2(n2802), .B0(ssrms0_out[23]), 
        .Y(pe_out[0]) );
  INVX2TS U3732 ( .A(reg_acc), .Y(n3146) );
  NOR2XLTS U3733 ( .A(n4789), .B(n3146), .Y(m1_out[0]) );
  NOR2XLTS U3734 ( .A(n4795), .B(n3146), .Y(m1_out[20]) );
  NOR2XLTS U3735 ( .A(n4794), .B(n3146), .Y(m1_out[3]) );
  NOR2XLTS U3736 ( .A(n4800), .B(n3146), .Y(m1_out[21]) );
  NOR2XLTS U3737 ( .A(n4799), .B(n3146), .Y(m1_out[1]) );
  NOR2XLTS U3738 ( .A(n4790), .B(n3146), .Y(m1_out[22]) );
  NOR2XLTS U3739 ( .A(n4804), .B(n3146), .Y(m1_out[2]) );
  NOR2XLTS U3740 ( .A(n4803), .B(n3146), .Y(m1_out[6]) );
  NOR2XLTS U3741 ( .A(n4802), .B(n3146), .Y(m1_out[10]) );
  NOR2XLTS U3742 ( .A(n4801), .B(n3146), .Y(m1_out[18]) );
  NOR2XLTS U3743 ( .A(n4788), .B(n3146), .Y(m1_out[12]) );
  NOR2XLTS U3744 ( .A(n4796), .B(n3146), .Y(m1_out[17]) );
  NOR2XLTS U3745 ( .A(n4797), .B(n3146), .Y(m1_out[13]) );
  NOR2XLTS U3746 ( .A(n4792), .B(n3146), .Y(m1_out[11]) );
  NOR2XLTS U3747 ( .A(n4793), .B(n3146), .Y(m1_out[7]) );
  NOR2XLTS U3748 ( .A(n4791), .B(n3146), .Y(m1_out[15]) );
  NOR2XLTS U3749 ( .A(n4798), .B(n3146), .Y(m1_out[5]) );
  NAND2X1TS U3750 ( .A(regindex_out[2]), .B(n3155), .Y(n3154) );
  NOR2XLTS U3751 ( .A(n4773), .B(n3154), .Y(n2805) );
  INVX2TS U3752 ( .A(mux13[0]), .Y(n4743) );
  NAND3XLTS U3753 ( .A(mux13[1]), .B(mux13[2]), .C(n4743), .Y(n3157) );
  AOI211XLTS U3754 ( .A0(n4773), .A1(n3154), .B0(n2805), .C0(n3157), .Y(
        m13_out[3]) );
  INVX2TS U3755 ( .A(n2805), .Y(n2807) );
  NAND2X1TS U3756 ( .A(regindex_out[4]), .B(n2805), .Y(n3158) );
  INVX2TS U3757 ( .A(n3158), .Y(n2806) );
  AOI211XLTS U3758 ( .A0(n4784), .A1(n2807), .B0(n2806), .C0(n3157), .Y(
        m13_out[4]) );
  CLKAND2X2TS U3759 ( .A(mux13[2]), .B(n4743), .Y(n2808) );
  INVX2TS U3760 ( .A(mux13[1]), .Y(n3153) );
  AO22XLTS U3761 ( .A0(n2809), .A1(n2808), .B0(mux13[2]), .B1(n3153), .Y(
        m13_out[1]) );
  INVX2TS U3762 ( .A(counterii[2]), .Y(n2810) );
  NAND2X1TS U3763 ( .A(counterii[1]), .B(n2810), .Y(n3799) );
  OAI21XLTS U3764 ( .A0(counterii[1]), .A1(n2810), .B0(n3799), .Y(n3798) );
  OA22X1TS U3765 ( .A0(\C43/DATA3_4 ), .A1(n3799), .B0(count_out[4]), .B1(
        n3798), .Y(n4779) );
  INVX2TS U3766 ( .A(sr_mp[0]), .Y(n3757) );
  NOR2XLTS U3767 ( .A(sr_mp[1]), .B(n3757), .Y(n2811) );
  BUFX3TS U3768 ( .A(n2811), .Y(n4413) );
  OR2X1TS U3769 ( .A(sr_mp[1]), .B(sr_mp[0]), .Y(n4304) );
  NAND2X1TS U3770 ( .A(sr_mp[1]), .B(sr_mp[0]), .Y(n3764) );
  AOI222XLTS U3771 ( .A0(n4413), .A1(mult2_out[0]), .B0(n1985), .B1(
        srmp_out[0]), .C0(n4412), .C1(srmp_out[1]), .Y(n2812) );
  INVX2TS U3772 ( .A(n2812), .Y(n1815) );
  AOI22X1TS U3773 ( .A0(n2316), .A1(n2819), .B0(n2816), .B1(n2818), .Y(n2832)
         );
  OAI22X1TS U3774 ( .A0(n2815), .A1(n2826), .B0(n3748), .B1(n2814), .Y(n2821)
         );
  INVX2TS U3775 ( .A(n2816), .Y(n2817) );
  OAI22X1TS U3776 ( .A0(n3739), .A1(n2819), .B0(n2818), .B1(n2817), .Y(n2820)
         );
  OAI32X1TS U3777 ( .A0(n2821), .A1(n3354), .A2(n2820), .B0(n2831), .B1(n2821), 
        .Y(n2830) );
  INVX2TS U3778 ( .A(n2822), .Y(n2824) );
  AOI21X1TS U3779 ( .A0(n2824), .A1(n2823), .B0(n3741), .Y(n2828) );
  OAI31X1TS U3780 ( .A0(n3728), .A1(n2828), .A2(n2827), .B0(n2826), .Y(n2829)
         );
  AOI22X1TS U3781 ( .A0(n2850), .A1(n3365), .B0(n2851), .B1(n2835), .Y(n2848)
         );
  NOR2BX1TS U3782 ( .AN(n2837), .B(n2836), .Y(n2845) );
  INVX2TS U3783 ( .A(n2846), .Y(n2843) );
  NOR2BX1TS U3784 ( .AN(n2839), .B(n2838), .Y(n2842) );
  OAI22X1TS U3785 ( .A0(n2850), .A1(n3422), .B0(n2845), .B1(n3741), .Y(n2840)
         );
  OAI32X1TS U3786 ( .A0(n2843), .A1(n2842), .A2(n3739), .B0(n2846), .B1(n2841), 
        .Y(n2844) );
  INVX2TS U3787 ( .A(n2858), .Y(n2853) );
  OAI32X1TS U3788 ( .A0(n2853), .A1(n2852), .A2(n2851), .B0(n3397), .B1(n2858), 
        .Y(n2867) );
  OAI2BB2XLTS U3789 ( .B0(n3741), .B1(n2859), .A0N(n2861), .A1N(n2316), .Y(
        n2864) );
  AOI22X1TS U3790 ( .A0(n3419), .A1(n2859), .B0(n3355), .B1(n2858), .Y(n2860)
         );
  INVX2TS U3791 ( .A(n2865), .Y(n2862) );
  AOI22X1TS U3792 ( .A0(n2865), .A1(n2864), .B0(n2863), .B1(n2862), .Y(n2866)
         );
  NOR2BX1TS U3793 ( .AN(n2870), .B(n2869), .Y(n2876) );
  NOR2BX1TS U3794 ( .AN(n2872), .B(n2871), .Y(n2874) );
  INVX2TS U3795 ( .A(n2455), .Y(n4714) );
  OAI22X1TS U3796 ( .A0(n2878), .A1(n4660), .B0(m17_out[1]), .B1(n4714), .Y(
        n2873) );
  AOI21X1TS U3797 ( .A0(n3526), .A1(m17_out[1]), .B0(n2873), .Y(n2880) );
  INVX2TS U3798 ( .A(n3503), .Y(n3306) );
  AOI22X1TS U3799 ( .A0(n2874), .A1(n3499), .B0(n3306), .B1(m17_out[1]), .Y(
        n2875) );
  AOI22X1TS U3800 ( .A0(n3493), .A1(n2878), .B0(m18_out[1]), .B1(n2877), .Y(
        n2879) );
  OAI32X1TS U3801 ( .A0(n2890), .A1(n2947), .A2(n2948), .B0(n2885), .B1(n2884), 
        .Y(n2899) );
  OAI2BB2XLTS U3802 ( .B0(n3741), .B1(n2891), .A0N(n2893), .A1N(n2316), .Y(
        n2896) );
  AOI22X1TS U3803 ( .A0(n3419), .A1(n2891), .B0(n3355), .B1(n2890), .Y(n2892)
         );
  INVX2TS U3804 ( .A(n2897), .Y(n2894) );
  AOI22X1TS U3805 ( .A0(n2897), .A1(n2896), .B0(n2895), .B1(n2894), .Y(n2898)
         );
  AOI22X1TS U3806 ( .A0(n3104), .A1(regep_out[8]), .B0(n3106), .B1(
        regeq_out[8]), .Y(n4717) );
  INVX2TS U3807 ( .A(n4717), .Y(m17_out[8]) );
  OAI32X1TS U3808 ( .A0(n2907), .A1(n2947), .A2(n2948), .B0(n2902), .B1(n2901), 
        .Y(n2916) );
  OAI2BB2XLTS U3809 ( .B0(n3741), .B1(n2908), .A0N(n2910), .A1N(n2316), .Y(
        n2913) );
  AOI22X1TS U3810 ( .A0(n3419), .A1(n2908), .B0(n3355), .B1(n2907), .Y(n2909)
         );
  INVX2TS U3811 ( .A(n2914), .Y(n2911) );
  AOI22X1TS U3812 ( .A0(n2914), .A1(n2913), .B0(n2912), .B1(n2911), .Y(n2915)
         );
  AOI22X1TS U3813 ( .A0(n3104), .A1(regep_out[10]), .B0(n3106), .B1(
        regeq_out[10]), .Y(n3486) );
  INVX2TS U3814 ( .A(n3486), .Y(m17_out[10]) );
  AOI22X1TS U3815 ( .A0(n3104), .A1(regep_out[20]), .B0(n3106), .B1(
        regeq_out[20]), .Y(n3608) );
  INVX2TS U3816 ( .A(n3608), .Y(m17_out[20]) );
  AOI22X1TS U3817 ( .A0(n3104), .A1(regep_out[19]), .B0(n3106), .B1(
        regeq_out[19]), .Y(n3120) );
  AOI22X1TS U3818 ( .A0(n3104), .A1(regep_out[18]), .B0(n3106), .B1(
        regeq_out[18]), .Y(n3574) );
  INVX2TS U3819 ( .A(n3574), .Y(m17_out[18]) );
  AOI22X1TS U3820 ( .A0(n3104), .A1(regep_out[16]), .B0(n3106), .B1(
        regeq_out[16]), .Y(n3541) );
  AOI22X1TS U3821 ( .A0(n3104), .A1(regep_out[17]), .B0(n3106), .B1(
        regeq_out[17]), .Y(n4691) );
  AOI22X1TS U3822 ( .A0(n3104), .A1(regep_out[15]), .B0(n3106), .B1(
        regeq_out[15]), .Y(n3552) );
  INVX2TS U3823 ( .A(n3552), .Y(m17_out[15]) );
  AOI22X1TS U3824 ( .A0(n3104), .A1(regep_out[14]), .B0(n3106), .B1(
        regeq_out[14]), .Y(n3560) );
  AOI22X1TS U3825 ( .A0(n3104), .A1(regep_out[13]), .B0(n3106), .B1(
        regeq_out[13]), .Y(n4703) );
  INVX2TS U3826 ( .A(n4703), .Y(m17_out[13]) );
  AOI22X1TS U3827 ( .A0(n3104), .A1(regep_out[12]), .B0(n3106), .B1(
        regeq_out[12]), .Y(n2938) );
  AOI22X1TS U3828 ( .A0(n3104), .A1(regep_out[11]), .B0(n3106), .B1(
        regeq_out[11]), .Y(n3523) );
  INVX2TS U3829 ( .A(n3523), .Y(m17_out[11]) );
  AOI22X1TS U3830 ( .A0(n3104), .A1(regep_out[9]), .B0(n3106), .B1(
        regeq_out[9]), .Y(n4721) );
  INVX2TS U3831 ( .A(n4721), .Y(m17_out[9]) );
  NAND2X1TS U3832 ( .A(n4717), .B(n3472), .Y(n4709) );
  NAND2X1TS U3833 ( .A(n3486), .B(n3482), .Y(n3520) );
  NAND2X1TS U3834 ( .A(n2938), .B(n3528), .Y(n4704) );
  NAND2X1TS U3835 ( .A(n3560), .B(n3557), .Y(n3565) );
  NAND2X1TS U3836 ( .A(n3120), .B(n2940), .Y(n3589) );
  NAND2X1TS U3837 ( .A(m17_out[9]), .B(n2925), .Y(n2924) );
  NAND2X1TS U3838 ( .A(n3547), .B(n2927), .Y(n2919) );
  INVX2TS U3839 ( .A(n2919), .Y(n2929) );
  INVX2TS U3840 ( .A(n3560), .Y(m17_out[14]) );
  INVX2TS U3841 ( .A(n4691), .Y(m17_out[17]) );
  NAND2X1TS U3842 ( .A(n2933), .B(m17_out[17]), .Y(n2932) );
  AOI21X1TS U3843 ( .A0(n3574), .A1(n2932), .B0(n2934), .Y(n3570) );
  AOI21X1TS U3844 ( .A0(n3541), .A1(n2930), .B0(n2933), .Y(n3538) );
  NAND2X1TS U3845 ( .A(n2929), .B(m17_out[13]), .Y(n2928) );
  NAND2X1TS U3846 ( .A(m17_out[13]), .B(m17_out[14]), .Y(n3550) );
  AOI21X1TS U3847 ( .A0(n3560), .A1(n2928), .B0(n2931), .Y(n3562) );
  NAND2X1TS U3848 ( .A(n2927), .B(m17_out[11]), .Y(n2926) );
  AOI21X1TS U3849 ( .A0(n2938), .A1(n2926), .B0(n2929), .Y(n3531) );
  AOI21X1TS U3850 ( .A0(n3486), .A1(n2924), .B0(n2927), .Y(n3487) );
  AOI21X1TS U3851 ( .A0(n4717), .A1(n2920), .B0(n2925), .Y(n3471) );
  NAND2X1TS U3852 ( .A(n4713), .B(n4712), .Y(n4711) );
  NAND2X1TS U3853 ( .A(n3518), .B(n3517), .Y(n3530) );
  NAND2X1TS U3854 ( .A(n4699), .B(n4698), .Y(n4697) );
  NAND2X1TS U3855 ( .A(n3561), .B(n3546), .Y(n3545) );
  NAND2X1TS U3856 ( .A(n4685), .B(n4684), .Y(n4683) );
  INVX2TS U3857 ( .A(n3120), .Y(m17_out[19]) );
  NAND2X1TS U3858 ( .A(n2934), .B(m17_out[19]), .Y(n3108) );
  NAND2X1TS U3859 ( .A(n3569), .B(n2935), .Y(n3583) );
  OAI32X1TS U3860 ( .A0(n2456), .A1(n3569), .A2(n2935), .B0(n3583), .B1(n2456), 
        .Y(n2945) );
  AOI21X1TS U3861 ( .A0(m18_out[7]), .A1(n2937), .B0(n2936), .Y(n4716) );
  NAND2X1TS U3862 ( .A(n4708), .B(m17_out[9]), .Y(n3483) );
  INVX2TS U3863 ( .A(n2938), .Y(m17_out[12]) );
  INVX2TS U3864 ( .A(n3541), .Y(m17_out[16]) );
  NAND2X1TS U3865 ( .A(n4688), .B(m17_out[16]), .Y(n4686) );
  NAND2X1TS U3866 ( .A(n3585), .B(m17_out[18]), .Y(n3119) );
  AOI21X1TS U3867 ( .A0(n4689), .A1(n3119), .B0(n2941), .Y(n2942) );
  AOI32X1TS U3868 ( .A0(n4714), .A1(n3120), .A2(n2943), .B0(n2942), .B1(
        m17_out[19]), .Y(n2944) );
  OR3X1TS U3869 ( .A(n2946), .B(n2945), .C(n2944), .Y(alutwo_out[19]) );
  AOI22X1TS U3870 ( .A0(n2950), .A1(n2968), .B0(n2997), .B1(n2998), .Y(n2963)
         );
  OAI2BB2XLTS U3871 ( .B0(n3741), .B1(n2955), .A0N(n2957), .A1N(n2316), .Y(
        n2960) );
  AOI22X1TS U3872 ( .A0(n3419), .A1(n2955), .B0(n3736), .B1(n2998), .Y(n2956)
         );
  INVX2TS U3873 ( .A(n2961), .Y(n2958) );
  AOI22X1TS U3874 ( .A0(n2961), .A1(n2960), .B0(n2959), .B1(n2958), .Y(n2962)
         );
  AOI22X1TS U3875 ( .A0(n2969), .A1(n2968), .B0(n2967), .B1(n2974), .Y(n2983)
         );
  OAI2BB2XLTS U3876 ( .B0(n3741), .B1(n2975), .A0N(n2977), .A1N(n2316), .Y(
        n2980) );
  AOI22X1TS U3877 ( .A0(n3419), .A1(n2975), .B0(n3355), .B1(n2974), .Y(n2976)
         );
  AOI22X1TS U3878 ( .A0(n2981), .A1(n2980), .B0(n2979), .B1(n2978), .Y(n2982)
         );
  AOI22X1TS U3879 ( .A0(n3104), .A1(regep_out[22]), .B0(n3106), .B1(
        regeq_out[22]), .Y(n3619) );
  INVX2TS U3880 ( .A(n3619), .Y(m17_out[22]) );
  AOI22X1TS U3881 ( .A0(n3104), .A1(regep_out[23]), .B0(n3106), .B1(
        regeq_out[23]), .Y(n4676) );
  INVX2TS U3882 ( .A(n4676), .Y(m17_out[23]) );
  AOI22X1TS U3883 ( .A0(n3104), .A1(regep_out[24]), .B0(n3106), .B1(
        regeq_out[24]), .Y(n4679) );
  INVX2TS U3884 ( .A(n4679), .Y(m17_out[24]) );
  NOR2BX1TS U3885 ( .AN(n2988), .B(n2987), .Y(n2990) );
  OAI22X1TS U3886 ( .A0(n2990), .A1(n3741), .B0(n3739), .B1(n2989), .Y(n2991)
         );
  OAI22X1TS U3887 ( .A0(n2996), .A1(n2993), .B0(n2992), .B1(n3748), .Y(n2994)
         );
  AOI21X1TS U3888 ( .A0(n2996), .A1(n2995), .B0(n2994), .Y(n3000) );
  AOI32X1TS U3889 ( .A0(n3729), .A1(n3001), .A2(n2998), .B0(n2997), .B1(n3001), 
        .Y(n2999) );
  NAND2X1TS U3890 ( .A(n3083), .B(n3003), .Y(n3024) );
  AOI22X1TS U3891 ( .A0(n3007), .A1(n3024), .B0(n3006), .B1(n3012), .Y(n3021)
         );
  OAI2BB2XLTS U3892 ( .B0(n3741), .B1(n3013), .A0N(n3015), .A1N(n2316), .Y(
        n3018) );
  AOI22X1TS U3893 ( .A0(n3419), .A1(n3013), .B0(n3736), .B1(n3012), .Y(n3014)
         );
  AOI22X1TS U3894 ( .A0(n3019), .A1(n3018), .B0(n3017), .B1(n3016), .Y(n3020)
         );
  AOI22X1TS U3895 ( .A0(n3104), .A1(regep_out[28]), .B0(n3106), .B1(
        regeq_out[28]), .Y(n3670) );
  INVX2TS U3896 ( .A(n3670), .Y(m17_out[28]) );
  AOI22X1TS U3897 ( .A0(n3104), .A1(regep_out[26]), .B0(n3106), .B1(
        regeq_out[26]), .Y(n3649) );
  INVX2TS U3898 ( .A(n3649), .Y(m17_out[26]) );
  AOI22X1TS U3899 ( .A0(n3104), .A1(regep_out[27]), .B0(n3106), .B1(
        regeq_out[27]), .Y(n3666) );
  INVX2TS U3900 ( .A(n3666), .Y(m17_out[27]) );
  AOI22X1TS U3901 ( .A0(n3025), .A1(n3024), .B0(n3023), .B1(n3030), .Y(n3039)
         );
  OAI2BB2XLTS U3902 ( .B0(n3741), .B1(n3031), .A0N(n3033), .A1N(n2316), .Y(
        n3036) );
  AOI22X1TS U3903 ( .A0(n3419), .A1(n3031), .B0(n3355), .B1(n3030), .Y(n3032)
         );
  AOI22X1TS U3904 ( .A0(n3037), .A1(n3036), .B0(n3035), .B1(n3034), .Y(n3038)
         );
  OAI2BB1X1TS U3905 ( .A0N(n3042), .A1N(n3041), .B0(n3083), .Y(n3063) );
  AOI22X1TS U3906 ( .A0(n3046), .A1(n3063), .B0(n3045), .B1(n3051), .Y(n3060)
         );
  OAI2BB2XLTS U3907 ( .B0(n3741), .B1(n3052), .A0N(n3054), .A1N(n2316), .Y(
        n3057) );
  AOI22X1TS U3908 ( .A0(n3419), .A1(n3052), .B0(n3736), .B1(n3051), .Y(n3053)
         );
  AOI22X1TS U3909 ( .A0(n3058), .A1(n3057), .B0(n3056), .B1(n3055), .Y(n3059)
         );
  AOI22X1TS U3910 ( .A0(n3064), .A1(n3063), .B0(n3062), .B1(n3069), .Y(n3078)
         );
  OAI2BB2XLTS U3911 ( .B0(n3741), .B1(n3070), .A0N(n3072), .A1N(n2316), .Y(
        n3075) );
  AOI22X1TS U3912 ( .A0(n3419), .A1(n3070), .B0(n3736), .B1(n3069), .Y(n3071)
         );
  AOI22X1TS U3913 ( .A0(n3076), .A1(n3075), .B0(n3074), .B1(n3073), .Y(n3077)
         );
  AOI22X1TS U3914 ( .A0(n3124), .A1(reges0_out[30]), .B0(n3125), .B1(
        srmt_out[30]), .Y(n3081) );
  AOI22X1TS U3915 ( .A0(n3123), .A1(regms_out[30]), .B0(n3122), .B1(
        regres_out[30]), .Y(n3080) );
  NAND2X1TS U3916 ( .A(n3081), .B(n3080), .Y(n3094) );
  INVX2TS U3917 ( .A(n3094), .Y(n3128) );
  AOI22X1TS U3918 ( .A0(n3128), .A1(n3732), .B0(n3086), .B1(n3094), .Y(n3102)
         );
  AOI222X1TS U3919 ( .A0(n2388), .A1(regms_out[30]), .B0(n2630), .B1(
        ssrms0_out[30]), .C0(n3132), .C1(srmt_out[30]), .Y(n3137) );
  OAI21XLTS U3920 ( .A0(n3092), .A1(n3088), .B0(n3087), .Y(n3089) );
  NAND2X1TS U3921 ( .A(n3094), .B(n3089), .Y(n3131) );
  AOI21X1TS U3922 ( .A0(n3092), .A1(n3091), .B0(n3090), .Y(n3093) );
  NAND2X1TS U3923 ( .A(n3093), .B(n3103), .Y(n3136) );
  OAI2BB2XLTS U3924 ( .B0(n3741), .B1(n3095), .A0N(n3097), .A1N(n2316), .Y(
        n3100) );
  AOI22X1TS U3925 ( .A0(n3419), .A1(n3095), .B0(n3736), .B1(n3094), .Y(n3096)
         );
  INVX2TS U3926 ( .A(n3137), .Y(n3098) );
  AOI22X1TS U3927 ( .A0(n3137), .A1(n3100), .B0(n3099), .B1(n3098), .Y(n3101)
         );
  CLKBUFX2TS U3928 ( .A(regmb_out[11]), .Y(n4815) );
  AO22XLTS U3929 ( .A0(n4612), .A1(regmc_out[1]), .B0(n4610), .B1(regma_out[1]), .Y(m19_out[1]) );
  AO22XLTS U3930 ( .A0(n4612), .A1(regmc_out[2]), .B0(n4610), .B1(regma_out[2]), .Y(m19_out[2]) );
  AO22XLTS U3931 ( .A0(n4612), .A1(regmc_out[3]), .B0(n4610), .B1(regma_out[3]), .Y(m19_out[3]) );
  AO22XLTS U3932 ( .A0(n4612), .A1(regmc_out[4]), .B0(n4610), .B1(regma_out[4]), .Y(m19_out[4]) );
  AO22XLTS U3933 ( .A0(n4612), .A1(regmc_out[5]), .B0(n4610), .B1(regma_out[5]), .Y(m19_out[5]) );
  AO22XLTS U3934 ( .A0(n4612), .A1(regmc_out[6]), .B0(n4610), .B1(regma_out[6]), .Y(m19_out[6]) );
  AO22XLTS U3935 ( .A0(n4612), .A1(regmc_out[7]), .B0(n4610), .B1(regma_out[7]), .Y(m19_out[7]) );
  AO22XLTS U3936 ( .A0(n4612), .A1(regmc_out[8]), .B0(n4610), .B1(regma_out[8]), .Y(m19_out[8]) );
  AO22XLTS U3937 ( .A0(n4612), .A1(regmc_out[9]), .B0(n4610), .B1(regma_out[9]), .Y(m19_out[9]) );
  AO22XLTS U3938 ( .A0(n4612), .A1(regmc_out[10]), .B0(n4610), .B1(
        regma_out[10]), .Y(m19_out[10]) );
  AO22XLTS U3939 ( .A0(n4612), .A1(regmc_out[11]), .B0(n4610), .B1(
        regma_out[11]), .Y(m19_out[11]) );
  AO22XLTS U3940 ( .A0(n4612), .A1(regmc_out[13]), .B0(n4610), .B1(
        regma_out[13]), .Y(m19_out[13]) );
  AO22XLTS U3941 ( .A0(n4612), .A1(regmc_out[14]), .B0(n4610), .B1(
        regma_out[14]), .Y(m19_out[14]) );
  CLKBUFX3TS U3942 ( .A(regmb_out[2]), .Y(n4814) );
  CLKBUFX2TS U3943 ( .A(regmb_out[17]), .Y(n4816) );
  AOI22X1TS U3944 ( .A0(n3104), .A1(regep_out[31]), .B0(n3106), .B1(
        regeq_out[31]), .Y(n3693) );
  INVX2TS U3945 ( .A(n3693), .Y(m17_out[31]) );
  AOI22X1TS U3946 ( .A0(n3104), .A1(regep_out[30]), .B0(n3106), .B1(
        regeq_out[30]), .Y(n4663) );
  INVX2TS U3947 ( .A(n4663), .Y(m17_out[30]) );
  AOI22X1TS U3948 ( .A0(n3104), .A1(regep_out[25]), .B0(n3106), .B1(
        regeq_out[25]), .Y(n3630) );
  INVX2TS U3949 ( .A(n3630), .Y(m17_out[25]) );
  NAND2X1TS U3950 ( .A(n3664), .B(m17_out[28]), .Y(n3105) );
  AOI22X1TS U3951 ( .A0(n3104), .A1(regep_out[21]), .B0(n3106), .B1(
        regeq_out[21]), .Y(n3611) );
  INVX2TS U3952 ( .A(n3611), .Y(m17_out[21]) );
  NAND2X1TS U3953 ( .A(n3110), .B(m17_out[21]), .Y(n3109) );
  NAND2X1TS U3954 ( .A(n3111), .B(m17_out[23]), .Y(n3112) );
  AOI22X1TS U3955 ( .A0(n3104), .A1(regep_out[29]), .B0(n3106), .B1(
        regeq_out[29]), .Y(n3680) );
  INVX2TS U3956 ( .A(n3680), .Y(m17_out[29]) );
  NAND2X1TS U3957 ( .A(n3118), .B(m17_out[29]), .Y(n3117) );
  AOI21X1TS U3958 ( .A0(n4663), .A1(n3117), .B0(n3690), .Y(n4667) );
  INVX2TS U3959 ( .A(n3112), .Y(n3107) );
  NAND2X1TS U3960 ( .A(n3664), .B(n3107), .Y(n3115) );
  AOI21X1TS U3961 ( .A0(n3670), .A1(n3115), .B0(n3118), .Y(n3662) );
  AOI21X1TS U3962 ( .A0(n3649), .A1(n3113), .B0(n3116), .Y(n3637) );
  AOI22X1TS U3963 ( .A0(n4679), .A1(n3112), .B0(n3107), .B1(m17_out[24]), .Y(
        n4672) );
  AOI21X1TS U3964 ( .A0(n3619), .A1(n3109), .B0(n3111), .Y(n3606) );
  AOI21X1TS U3965 ( .A0(n3608), .A1(n3108), .B0(n3110), .Y(n3584) );
  NAND2X1TS U3966 ( .A(n3597), .B(n3596), .Y(n3605) );
  NAND2X1TS U3967 ( .A(n3621), .B(n3620), .Y(n4671) );
  NAND2X1TS U3968 ( .A(n4670), .B(n3626), .Y(n3636) );
  NAND2X1TS U3969 ( .A(n3647), .B(n3646), .Y(n3661) );
  NAND2X1TS U3970 ( .A(n3678), .B(n3677), .Y(n3676) );
  NAND2X1TS U3971 ( .A(n3611), .B(n3593), .Y(n3609) );
  NAND2X1TS U3972 ( .A(n4710), .B(n3622), .Y(n3639) );
  NAND2X1TS U3973 ( .A(n3670), .B(n3671), .Y(n3686) );
  NAND2X1TS U3974 ( .A(n4663), .B(n4661), .Y(n3697) );
  AOI21X1TS U3975 ( .A0(n4696), .A1(n3692), .B0(n3695), .Y(n4669) );
  NOR2BX1TS U3976 ( .AN(n3676), .B(n2456), .Y(n4666) );
  NAND2X1TS U3977 ( .A(n3682), .B(m17_out[29]), .Y(n4664) );
  AOI32X1TS U3978 ( .A0(n3690), .A1(m17_out[31]), .A2(n4666), .B0(n3694), .B1(
        m17_out[31]), .Y(n3121) );
  OAI31X1TS U3979 ( .A0(n4669), .A1(m17_out[31]), .A2(m17_out[30]), .B0(n3121), 
        .Y(\alutwo/N325 ) );
  AOI22X1TS U3980 ( .A0(regms_out[31]), .A1(n3123), .B0(n3122), .B1(
        regres_out[31]), .Y(n3127) );
  AOI22X1TS U3981 ( .A0(srmt_out[31]), .A1(n3125), .B0(n3124), .B1(
        reges0_out[31]), .Y(n3126) );
  NAND2X1TS U3982 ( .A(n3127), .B(n3126), .Y(n3735) );
  INVX2TS U3983 ( .A(n3735), .Y(n3145) );
  INVX2TS U3984 ( .A(n3140), .Y(n3144) );
  AOI21X1TS U3985 ( .A0(n3137), .A1(n3131), .B0(n3130), .Y(n3734) );
  AOI222XLTS U3986 ( .A0(ssrms0_out[31]), .A1(n2630), .B0(regms_out[31]), .B1(
        n2388), .C0(srmt_out[31]), .C1(n3132), .Y(n3743) );
  INVX2TS U3987 ( .A(n3743), .Y(n3138) );
  AOI222XLTS U3988 ( .A0(n3734), .A1(n3735), .B0(n3734), .B1(n3138), .C0(n3735), .C1(n3138), .Y(n3134) );
  OAI32X1TS U3989 ( .A0(alu1[0]), .A1(n3735), .A2(n3730), .B0(n3134), .B1(
        n3133), .Y(n3142) );
  AOI21X1TS U3990 ( .A0(n3137), .A1(n3136), .B0(n3135), .Y(n3733) );
  AOI222XLTS U3991 ( .A0(n3733), .A1(n3138), .B0(n3733), .B1(n3749), .C0(n3138), .C1(n3749), .Y(n3139) );
  AOI211XLTS U3992 ( .A0(n3140), .A1(n3735), .B0(n3739), .C0(n3139), .Y(n3141)
         );
  AOI31XLTS U3993 ( .A0(\aluone/N324 ), .A1(n3142), .A2(n3424), .B0(n3141), 
        .Y(n3143) );
  OAI31X1TS U3994 ( .A0(n3145), .A1(n3144), .A2(n3748), .B0(n3143), .Y(
        \aluone/N325 ) );
  NOR2XLTS U3995 ( .A(n4786), .B(n3146), .Y(m1_out[29]) );
  NOR2XLTS U3996 ( .A(n4785), .B(n3146), .Y(m1_out[23]) );
  NOR2XLTS U3997 ( .A(n4775), .B(n3146), .Y(m1_out[24]) );
  NOR2XLTS U3998 ( .A(n4781), .B(n3146), .Y(m1_out[25]) );
  NOR2XLTS U3999 ( .A(n4782), .B(n3146), .Y(m1_out[26]) );
  NOR2XLTS U4000 ( .A(n4776), .B(n3146), .Y(m1_out[28]) );
  NOR2XLTS U4001 ( .A(n4783), .B(n3146), .Y(m1_out[30]) );
  INVX2TS U4002 ( .A(mux6[1]), .Y(n3148) );
  OAI21XLTS U4003 ( .A0(regss_out), .A1(n3148), .B0(mux6[0]), .Y(n3149) );
  OAI21XLTS U4004 ( .A0(regst_out), .A1(n3148), .B0(n3149), .Y(n3147) );
  OAI31X1TS U4005 ( .A0(regst_out), .A1(n3149), .A2(n3148), .B0(n3147), .Y(
        \m6_out[0] ) );
  NAND2X1TS U4006 ( .A(reg_i), .B(mux22), .Y(n4607) );
  OAI21XLTS U4007 ( .A0(reg_i), .A1(n4813), .B0(n4607), .Y(n1686) );
  AOI2BB1XLTS U4008 ( .A0N(regindex_out[0]), .A1N(regi_out[0]), .B0(n3150), 
        .Y(n3151) );
  OAI211XLTS U4009 ( .A0(n3151), .A1(n3153), .B0(mux13[2]), .C0(n4743), .Y(
        n3152) );
  OAI31X1TS U4010 ( .A0(mux13[2]), .A1(n4743), .A2(n3153), .B0(n3152), .Y(
        m13_out[0]) );
  OAI21XLTS U4011 ( .A0(regindex_out[2]), .A1(n3155), .B0(n3154), .Y(n3156) );
  NOR2XLTS U4012 ( .A(n3157), .B(n3156), .Y(m13_out[2]) );
  AOI211XLTS U4013 ( .A0(n4774), .A1(n3158), .B0(Coutadd), .C0(n3157), .Y(
        m13_out[5]) );
  NOR3X1TS U4014 ( .A(mux3[2]), .B(mux13[0]), .C(mux3[1]), .Y(n4739) );
  INVX1TS U4015 ( .A(n4739), .Y(n3159) );
  NOR3BX1TS U4016 ( .AN(mux3[2]), .B(mux13[0]), .C(mux3[1]), .Y(n3178) );
  NAND2BXLTS U4017 ( .AN(mux3[2]), .B(mux3[1]), .Y(n4741) );
  NOR2X2TS U4018 ( .A(mux13[0]), .B(n4741), .Y(n3411) );
  AOI22X1TS U4019 ( .A0(n3178), .A1(srmp_out[33]), .B0(n3411), .B1(rf_aout[10]), .Y(n3160) );
  OAI21XLTS U4020 ( .A0(n3159), .A1(n4802), .B0(n3160), .Y(m3_out[10]) );
  AOI22X1TS U4021 ( .A0(n3178), .A1(srmp_out[24]), .B0(n3411), .B1(rf_aout[1]), 
        .Y(n3161) );
  OAI21XLTS U4022 ( .A0(n3159), .A1(n4799), .B0(n3161), .Y(m3_out[1]) );
  AOI22X1TS U4023 ( .A0(n3178), .A1(srmp_out[28]), .B0(n3411), .B1(rf_aout[5]), 
        .Y(n3162) );
  OAI21XLTS U4024 ( .A0(n3159), .A1(n4798), .B0(n3162), .Y(m3_out[5]) );
  AOI22X1TS U4025 ( .A0(n3178), .A1(srmp_out[26]), .B0(n3411), .B1(rf_aout[3]), 
        .Y(n3163) );
  OAI21XLTS U4026 ( .A0(n3159), .A1(n4794), .B0(n3163), .Y(m3_out[3]) );
  INVX2TS U4027 ( .A(n3799), .Y(n4819) );
  AOI22X1TS U4028 ( .A0(n3178), .A1(srmp_out[30]), .B0(n3411), .B1(rf_aout[7]), 
        .Y(n3164) );
  OAI21XLTS U4029 ( .A0(n3159), .A1(n4793), .B0(n3164), .Y(m3_out[7]) );
  AOI22X1TS U4030 ( .A0(n3178), .A1(srmp_out[35]), .B0(n3411), .B1(rf_aout[12]), .Y(n3165) );
  OAI21XLTS U4031 ( .A0(n3159), .A1(n4788), .B0(n3165), .Y(m3_out[12]) );
  AOI22X1TS U4032 ( .A0(n3178), .A1(srmp_out[29]), .B0(n3411), .B1(rf_aout[6]), 
        .Y(n3166) );
  OAI21XLTS U4033 ( .A0(n3159), .A1(n4803), .B0(n3166), .Y(m3_out[6]) );
  AOI22X1TS U4034 ( .A0(n3178), .A1(srmp_out[25]), .B0(n3411), .B1(rf_aout[2]), 
        .Y(n3167) );
  OAI21XLTS U4035 ( .A0(n3159), .A1(n4804), .B0(n3167), .Y(m3_out[2]) );
  AOI22X1TS U4036 ( .A0(n3178), .A1(srmp_out[34]), .B0(n3411), .B1(rf_aout[11]), .Y(n3168) );
  OAI21XLTS U4037 ( .A0(n3159), .A1(n4792), .B0(n3168), .Y(m3_out[11]) );
  INVX2TS U4038 ( .A(mux2[1]), .Y(n4725) );
  INVX2TS U4039 ( .A(mux2[2]), .Y(n3174) );
  NAND2X1TS U4040 ( .A(n4725), .B(n3174), .Y(n3230) );
  NOR3X1TS U4041 ( .A(mux2[0]), .B(n4725), .C(n3174), .Y(n3259) );
  CLKBUFX2TS U4042 ( .A(n3259), .Y(n4731) );
  NAND2X1TS U4043 ( .A(mux2[0]), .B(n3174), .Y(n3231) );
  INVX2TS U4044 ( .A(rf_aout[26]), .Y(n3444) );
  INVX2TS U4045 ( .A(mux2[0]), .Y(n3218) );
  NAND3XLTS U4046 ( .A(mux2[2]), .B(n4725), .C(n3218), .Y(n3264) );
  OAI22X1TS U4047 ( .A0(n3169), .A1(n3231), .B0(n3444), .B1(n3264), .Y(n3170)
         );
  AOI21X1TS U4048 ( .A0(n4731), .A1(regreg_out[26]), .B0(n3170), .Y(n3172) );
  NOR2X1TS U4049 ( .A(n3218), .B(mux2[1]), .Y(n4729) );
  OAI21XLTS U4050 ( .A0(regacc_out[26]), .A1(n3174), .B0(n4729), .Y(n3171) );
  OAI211XLTS U4051 ( .A0(n3230), .A1(n4806), .B0(n3172), .C0(n3171), .Y(
        m2_out[26]) );
  INVX2TS U4052 ( .A(ssrms0_out[11]), .Y(n4204) );
  NOR2X1TS U4053 ( .A(n4725), .B(n3231), .Y(n3260) );
  INVX2TS U4054 ( .A(n3260), .Y(n3258) );
  OR2X1TS U4055 ( .A(mux2[0]), .B(n3230), .Y(n3173) );
  INVX2TS U4056 ( .A(n3173), .Y(n3261) );
  AOI22X1TS U4057 ( .A0(n3259), .A1(regreg_out[11]), .B0(n3261), .B1(
        regcurrterm_out[11]), .Y(n3177) );
  INVX2TS U4058 ( .A(n3264), .Y(n4732) );
  AOI22X1TS U4059 ( .A0(n4732), .A1(rf_aout[11]), .B0(n3175), .B1(
        regacc_out[11]), .Y(n3176) );
  OAI211XLTS U4060 ( .A0(n4204), .A1(n3258), .B0(n3177), .C0(n3176), .Y(
        m2_out[11]) );
  INVX2TS U4061 ( .A(n3411), .Y(n3193) );
  INVX2TS U4062 ( .A(rf_aout[8]), .Y(n3290) );
  CLKBUFX2TS U4063 ( .A(n3178), .Y(n4740) );
  AOI22X1TS U4064 ( .A0(n4740), .A1(srmp_out[31]), .B0(n4739), .B1(
        regsum_out[8]), .Y(n3179) );
  OAI21XLTS U4065 ( .A0(n3193), .A1(n3290), .B0(n3179), .Y(m3_out[8]) );
  AOI22X1TS U4066 ( .A0(n4740), .A1(srmp_out[23]), .B0(n3411), .B1(rf_aout[0]), 
        .Y(n3180) );
  OAI21XLTS U4067 ( .A0(n3159), .A1(n4789), .B0(n3180), .Y(m3_out[0]) );
  INVX2TS U4068 ( .A(rf_aout[4]), .Y(n3296) );
  AOI22X1TS U4069 ( .A0(n4740), .A1(srmp_out[27]), .B0(n4739), .B1(
        regsum_out[4]), .Y(n3181) );
  OAI21XLTS U4070 ( .A0(n3193), .A1(n3296), .B0(n3181), .Y(m3_out[4]) );
  AOI22X1TS U4071 ( .A0(n4740), .A1(srmp_out[41]), .B0(n3411), .B1(rf_aout[18]), .Y(n3182) );
  OAI21XLTS U4072 ( .A0(n3159), .A1(n4801), .B0(n3182), .Y(m3_out[18]) );
  AOI22X1TS U4073 ( .A0(n4740), .A1(srmp_out[36]), .B0(n3411), .B1(rf_aout[13]), .Y(n3183) );
  OAI21XLTS U4074 ( .A0(n3159), .A1(n4797), .B0(n3183), .Y(m3_out[13]) );
  INVX2TS U4075 ( .A(rf_aout[14]), .Y(n3292) );
  AOI22X1TS U4076 ( .A0(n4740), .A1(srmp_out[37]), .B0(n4739), .B1(
        regsum_out[14]), .Y(n3184) );
  OAI21XLTS U4077 ( .A0(n3193), .A1(n3292), .B0(n3184), .Y(m3_out[14]) );
  INVX2TS U4078 ( .A(rf_aout[31]), .Y(n3237) );
  AOI22X1TS U4079 ( .A0(n4740), .A1(regsp_out), .B0(n4739), .B1(regsum_out[31]), .Y(n3185) );
  OAI21XLTS U4080 ( .A0(n3193), .A1(n3237), .B0(n3185), .Y(m3_out[31]) );
  INVX2TS U4081 ( .A(rf_aout[9]), .Y(n3288) );
  AOI22X1TS U4082 ( .A0(n4740), .A1(srmp_out[32]), .B0(n4739), .B1(
        regsum_out[9]), .Y(n3186) );
  OAI21XLTS U4083 ( .A0(n3193), .A1(n3288), .B0(n3186), .Y(m3_out[9]) );
  INVX2TS U4084 ( .A(rf_aout[16]), .Y(n3294) );
  AOI22X1TS U4085 ( .A0(n4740), .A1(srmp_out[39]), .B0(n4739), .B1(
        regsum_out[16]), .Y(n3187) );
  OAI21XLTS U4086 ( .A0(n3193), .A1(n3294), .B0(n3187), .Y(m3_out[16]) );
  AOI22X1TS U4087 ( .A0(n4740), .A1(srmp_out[40]), .B0(n3411), .B1(rf_aout[17]), .Y(n3188) );
  OAI21XLTS U4088 ( .A0(n3159), .A1(n4796), .B0(n3188), .Y(m3_out[17]) );
  AOI22X1TS U4089 ( .A0(n4740), .A1(srmp_out[45]), .B0(n3411), .B1(rf_aout[22]), .Y(n3189) );
  OAI21XLTS U4090 ( .A0(n3159), .A1(n4790), .B0(n3189), .Y(m3_out[22]) );
  AOI22X1TS U4091 ( .A0(n4740), .A1(srmp_out[44]), .B0(n3411), .B1(rf_aout[21]), .Y(n3190) );
  OAI21XLTS U4092 ( .A0(n3159), .A1(n4800), .B0(n3190), .Y(m3_out[21]) );
  AOI22X1TS U4093 ( .A0(n4740), .A1(srmp_out[43]), .B0(n3411), .B1(rf_aout[20]), .Y(n3191) );
  OAI21XLTS U4094 ( .A0(n3159), .A1(n4795), .B0(n3191), .Y(m3_out[20]) );
  INVX2TS U4095 ( .A(rf_aout[19]), .Y(n3298) );
  AOI22X1TS U4096 ( .A0(n4740), .A1(srmp_out[42]), .B0(n4739), .B1(
        regsum_out[19]), .Y(n3192) );
  OAI21XLTS U4097 ( .A0(n3193), .A1(n3298), .B0(n3192), .Y(m3_out[19]) );
  AOI22X1TS U4098 ( .A0(n4740), .A1(srmp_out[38]), .B0(n3411), .B1(rf_aout[15]), .Y(n3194) );
  OAI21XLTS U4099 ( .A0(n3159), .A1(n4791), .B0(n3194), .Y(m3_out[15]) );
  AOI22X1TS U4100 ( .A0(n4732), .A1(rf_aout[21]), .B0(n3175), .B1(
        regacc_out[21]), .Y(n3196) );
  AOI22X1TS U4101 ( .A0(n3259), .A1(regreg_out[21]), .B0(n3261), .B1(
        regcurrterm_out[21]), .Y(n3195) );
  OAI211XLTS U4102 ( .A0(n4100), .A1(n3258), .B0(n3196), .C0(n3195), .Y(
        m2_out[21]) );
  INVX2TS U4103 ( .A(ssrms0_out[1]), .Y(n4300) );
  AOI22X1TS U4104 ( .A0(n4732), .A1(rf_aout[1]), .B0(n3175), .B1(regacc_out[1]), .Y(n3198) );
  AOI22X1TS U4105 ( .A0(n3259), .A1(regreg_out[1]), .B0(n3261), .B1(
        regcurrterm_out[1]), .Y(n3197) );
  OAI211XLTS U4106 ( .A0(n4300), .A1(n3258), .B0(n3198), .C0(n3197), .Y(
        m2_out[1]) );
  AOI22X1TS U4107 ( .A0(n3175), .A1(regacc_out[2]), .B0(n3259), .B1(
        regreg_out[2]), .Y(n3200) );
  AOI22X1TS U4108 ( .A0(n4732), .A1(rf_aout[2]), .B0(n3261), .B1(
        regcurrterm_out[2]), .Y(n3199) );
  OAI211XLTS U4109 ( .A0(n4286), .A1(n3258), .B0(n3200), .C0(n3199), .Y(
        m2_out[2]) );
  AOI22X1TS U4110 ( .A0(n4732), .A1(rf_aout[7]), .B0(n3175), .B1(regacc_out[7]), .Y(n3202) );
  AOI22X1TS U4111 ( .A0(n3259), .A1(regreg_out[7]), .B0(n3261), .B1(
        regcurrterm_out[7]), .Y(n3201) );
  OAI211XLTS U4112 ( .A0(n4239), .A1(n3258), .B0(n3202), .C0(n3201), .Y(
        m2_out[7]) );
  AOI22X1TS U4113 ( .A0(n4732), .A1(rf_aout[12]), .B0(n3175), .B1(
        regacc_out[12]), .Y(n3204) );
  AOI22X1TS U4114 ( .A0(n3259), .A1(regreg_out[12]), .B0(n3261), .B1(
        regcurrterm_out[12]), .Y(n3203) );
  OAI211XLTS U4115 ( .A0(n4196), .A1(n3258), .B0(n3204), .C0(n3203), .Y(
        m2_out[12]) );
  INVX2TS U4116 ( .A(ssrms0_out[10]), .Y(n4213) );
  AOI22X1TS U4117 ( .A0(n3175), .A1(regacc_out[10]), .B0(n4731), .B1(
        regreg_out[10]), .Y(n3206) );
  AOI22X1TS U4118 ( .A0(n4732), .A1(rf_aout[10]), .B0(n3261), .B1(
        regcurrterm_out[10]), .Y(n3205) );
  OAI211XLTS U4119 ( .A0(n4213), .A1(n3258), .B0(n3206), .C0(n3205), .Y(
        m2_out[10]) );
  AOI22X1TS U4120 ( .A0(n3175), .A1(regacc_out[3]), .B0(n3259), .B1(
        regreg_out[3]), .Y(n3208) );
  AOI22X1TS U4121 ( .A0(n4732), .A1(rf_aout[3]), .B0(n3261), .B1(
        regcurrterm_out[3]), .Y(n3207) );
  OAI211XLTS U4122 ( .A0(n4276), .A1(n3258), .B0(n3208), .C0(n3207), .Y(
        m2_out[3]) );
  AOI22X1TS U4123 ( .A0(n4732), .A1(rf_aout[18]), .B0(n3175), .B1(
        regacc_out[18]), .Y(n3210) );
  AOI22X1TS U4124 ( .A0(n3259), .A1(regreg_out[18]), .B0(n3261), .B1(
        regcurrterm_out[18]), .Y(n3209) );
  OAI211XLTS U4125 ( .A0(n4137), .A1(n3258), .B0(n3210), .C0(n3209), .Y(
        m2_out[18]) );
  INVX2TS U4126 ( .A(ssrms0_out[0]), .Y(n3961) );
  AOI22X1TS U4127 ( .A0(n3175), .A1(regacc_out[0]), .B0(n4731), .B1(
        regreg_out[0]), .Y(n3212) );
  AOI22X1TS U4128 ( .A0(n4732), .A1(rf_aout[0]), .B0(n3261), .B1(
        regcurrterm_out[0]), .Y(n3211) );
  OAI211XLTS U4129 ( .A0(n3961), .A1(n3258), .B0(n3212), .C0(n3211), .Y(
        m2_out[0]) );
  INVX2TS U4130 ( .A(rf_aout[29]), .Y(n4737) );
  AOI21X1TS U4131 ( .A0(n4805), .A1(n3218), .B0(n3230), .Y(n3213) );
  AOI21X1TS U4132 ( .A0(regacc_out[29]), .A1(n4729), .B0(n3213), .Y(n3215) );
  INVX2TS U4133 ( .A(n3231), .Y(n4730) );
  AOI22X1TS U4134 ( .A0(reges0_out[6]), .A1(n4730), .B0(n4731), .B1(
        regreg_out[29]), .Y(n3214) );
  OAI211XLTS U4135 ( .A0(n4737), .A1(n3264), .B0(n3215), .C0(n3214), .Y(
        m2_out[29]) );
  AOI22X1TS U4136 ( .A0(n3175), .A1(regacc_out[13]), .B0(n3261), .B1(
        regcurrterm_out[13]), .Y(n3217) );
  AOI22X1TS U4137 ( .A0(n4732), .A1(rf_aout[13]), .B0(n4731), .B1(
        regreg_out[13]), .Y(n3216) );
  OAI211XLTS U4138 ( .A0(n4189), .A1(n3258), .B0(n3217), .C0(n3216), .Y(
        m2_out[13]) );
  INVX2TS U4139 ( .A(rf_aout[25]), .Y(n3416) );
  AOI21X1TS U4140 ( .A0(n4787), .A1(n3218), .B0(n3230), .Y(n3219) );
  AOI21X1TS U4141 ( .A0(regacc_out[25]), .A1(n4729), .B0(n3219), .Y(n3221) );
  AOI22X1TS U4142 ( .A0(reges0_out[2]), .A1(n4730), .B0(n4731), .B1(
        regreg_out[25]), .Y(n3220) );
  OAI211XLTS U4143 ( .A0(n3416), .A1(n3264), .B0(n3221), .C0(n3220), .Y(
        m2_out[25]) );
  INVX2TS U4144 ( .A(rf_aout[30]), .Y(n3513) );
  AOI22X1TS U4145 ( .A0(regcurrterm_out[30]), .A1(n3261), .B0(n3175), .B1(
        regacc_out[30]), .Y(n3223) );
  AOI22X1TS U4146 ( .A0(reges0_out[7]), .A1(n3260), .B0(n4731), .B1(
        regreg_out[30]), .Y(n3222) );
  OAI211XLTS U4147 ( .A0(n3513), .A1(n3264), .B0(n3223), .C0(n3222), .Y(
        m2_out[30]) );
  AOI2BB1XLTS U4148 ( .A0N(regcurrterm_out[28]), .A1N(mux2[0]), .B0(n3230), 
        .Y(n3224) );
  AOI21X1TS U4149 ( .A0(n4729), .A1(regacc_out[28]), .B0(n3224), .Y(n3226) );
  AOI22X1TS U4150 ( .A0(rf_aout[28]), .A1(n4732), .B0(n4731), .B1(
        regreg_out[28]), .Y(n3225) );
  OAI211XLTS U4151 ( .A0(n3227), .A1(n3231), .B0(n3226), .C0(n3225), .Y(
        m2_out[28]) );
  AOI22X1TS U4152 ( .A0(ssrms0_out[14]), .A1(n3260), .B0(n3261), .B1(
        regcurrterm_out[14]), .Y(n3229) );
  AOI22X1TS U4153 ( .A0(n3175), .A1(regacc_out[14]), .B0(n4731), .B1(
        regreg_out[14]), .Y(n3228) );
  OAI211XLTS U4154 ( .A0(n3264), .A1(n3292), .B0(n3229), .C0(n3228), .Y(
        m2_out[14]) );
  INVX2TS U4155 ( .A(rf_aout[23]), .Y(n3414) );
  INVX2TS U4156 ( .A(n3230), .Y(n4733) );
  AOI2BB1XLTS U4157 ( .A0N(n4725), .A1N(reges0_out[0]), .B0(n3231), .Y(n3232)
         );
  AOI21X1TS U4158 ( .A0(n4733), .A1(regcurrterm_out[23]), .B0(n3232), .Y(n3234) );
  AOI22X1TS U4159 ( .A0(n4729), .A1(regacc_out[23]), .B0(n4731), .B1(
        regreg_out[23]), .Y(n3233) );
  OAI211XLTS U4160 ( .A0(n3414), .A1(n3264), .B0(n3234), .C0(n3233), .Y(
        m2_out[23]) );
  AOI22X1TS U4161 ( .A0(n3260), .A1(regss0_out), .B0(n3261), .B1(
        regcurrterm_out[31]), .Y(n3236) );
  AOI22X1TS U4162 ( .A0(n3175), .A1(regacc_out[31]), .B0(n4731), .B1(
        regreg_out[31]), .Y(n3235) );
  OAI211XLTS U4163 ( .A0(n3237), .A1(n3264), .B0(n3236), .C0(n3235), .Y(
        m2_out[31]) );
  AOI22X1TS U4164 ( .A0(n4732), .A1(rf_aout[6]), .B0(n3261), .B1(
        regcurrterm_out[6]), .Y(n3239) );
  AOI22X1TS U4165 ( .A0(n3175), .A1(regacc_out[6]), .B0(n4731), .B1(
        regreg_out[6]), .Y(n3238) );
  OAI211XLTS U4166 ( .A0(n4248), .A1(n3258), .B0(n3239), .C0(n3238), .Y(
        m2_out[6]) );
  AOI22X1TS U4167 ( .A0(ssrms0_out[19]), .A1(n3260), .B0(n3261), .B1(
        regcurrterm_out[19]), .Y(n3241) );
  AOI22X1TS U4168 ( .A0(n3175), .A1(regacc_out[19]), .B0(n4731), .B1(
        regreg_out[19]), .Y(n3240) );
  OAI211XLTS U4169 ( .A0(n3264), .A1(n3298), .B0(n3241), .C0(n3240), .Y(
        m2_out[19]) );
  INVX2TS U4170 ( .A(ssrms0_out[22]), .Y(n4091) );
  AOI22X1TS U4171 ( .A0(n4732), .A1(rf_aout[22]), .B0(n3261), .B1(
        regcurrterm_out[22]), .Y(n3243) );
  AOI22X1TS U4172 ( .A0(n3175), .A1(regacc_out[22]), .B0(n4731), .B1(
        regreg_out[22]), .Y(n3242) );
  OAI211XLTS U4173 ( .A0(n4091), .A1(n3258), .B0(n3243), .C0(n3242), .Y(
        m2_out[22]) );
  AOI22X1TS U4174 ( .A0(n4732), .A1(rf_aout[17]), .B0(n3261), .B1(
        regcurrterm_out[17]), .Y(n3245) );
  AOI22X1TS U4175 ( .A0(n3175), .A1(regacc_out[17]), .B0(n4731), .B1(
        regreg_out[17]), .Y(n3244) );
  OAI211XLTS U4176 ( .A0(n4147), .A1(n3258), .B0(n3245), .C0(n3244), .Y(
        m2_out[17]) );
  AOI22X1TS U4177 ( .A0(ssrms0_out[9]), .A1(n3260), .B0(n3261), .B1(
        regcurrterm_out[9]), .Y(n3247) );
  AOI22X1TS U4178 ( .A0(n3175), .A1(regacc_out[9]), .B0(n4731), .B1(
        regreg_out[9]), .Y(n3246) );
  OAI211XLTS U4179 ( .A0(n3264), .A1(n3288), .B0(n3247), .C0(n3246), .Y(
        m2_out[9]) );
  AOI22X1TS U4180 ( .A0(ssrms0_out[4]), .A1(n3260), .B0(n3261), .B1(
        regcurrterm_out[4]), .Y(n3249) );
  AOI22X1TS U4181 ( .A0(n3175), .A1(regacc_out[4]), .B0(n4731), .B1(
        regreg_out[4]), .Y(n3248) );
  OAI211XLTS U4182 ( .A0(n3264), .A1(n3296), .B0(n3249), .C0(n3248), .Y(
        m2_out[4]) );
  AOI22X1TS U4183 ( .A0(n4732), .A1(rf_aout[5]), .B0(n3261), .B1(
        regcurrterm_out[5]), .Y(n3251) );
  AOI22X1TS U4184 ( .A0(n3175), .A1(regacc_out[5]), .B0(n4731), .B1(
        regreg_out[5]), .Y(n3250) );
  OAI211XLTS U4185 ( .A0(n4257), .A1(n3258), .B0(n3251), .C0(n3250), .Y(
        m2_out[5]) );
  AOI22X1TS U4186 ( .A0(ssrms0_out[16]), .A1(n3260), .B0(n3261), .B1(
        regcurrterm_out[16]), .Y(n3253) );
  AOI22X1TS U4187 ( .A0(n3175), .A1(regacc_out[16]), .B0(n4731), .B1(
        regreg_out[16]), .Y(n3252) );
  OAI211XLTS U4188 ( .A0(n3264), .A1(n3294), .B0(n3253), .C0(n3252), .Y(
        m2_out[16]) );
  AOI22X1TS U4189 ( .A0(ssrms0_out[20]), .A1(n3260), .B0(n4732), .B1(
        rf_aout[20]), .Y(n3255) );
  AOI22X1TS U4190 ( .A0(n3175), .A1(regacc_out[20]), .B0(n4731), .B1(
        regreg_out[20]), .Y(n3254) );
  OAI211XLTS U4191 ( .A0(n3173), .A1(n4807), .B0(n3255), .C0(n3254), .Y(
        m2_out[20]) );
  AOI22X1TS U4192 ( .A0(n4732), .A1(rf_aout[15]), .B0(n4731), .B1(
        regreg_out[15]), .Y(n3257) );
  AOI22X1TS U4193 ( .A0(n3175), .A1(regacc_out[15]), .B0(n3261), .B1(
        regcurrterm_out[15]), .Y(n3256) );
  OAI211XLTS U4194 ( .A0(n4175), .A1(n3258), .B0(n3257), .C0(n3256), .Y(
        m2_out[15]) );
  AOI22X1TS U4195 ( .A0(ssrms0_out[8]), .A1(n3260), .B0(n3259), .B1(
        regreg_out[8]), .Y(n3263) );
  AOI22X1TS U4196 ( .A0(n3175), .A1(regacc_out[8]), .B0(n3261), .B1(
        regcurrterm_out[8]), .Y(n3262) );
  OAI211XLTS U4197 ( .A0(n3264), .A1(n3290), .B0(n3263), .C0(n3262), .Y(
        m2_out[8]) );
  NAND2BXLTS U4198 ( .AN(ssr_ms0[1]), .B(ssr_ms0[0]), .Y(n3276) );
  NOR3BX1TS U4199 ( .AN(mux12[0]), .B(n3276), .C(mux12[1]), .Y(n4145) );
  NAND2X1TS U4200 ( .A(n4772), .B(n4778), .Y(n4082) );
  INVX2TS U4201 ( .A(n4082), .Y(n4160) );
  NAND2X1TS U4202 ( .A(n4145), .B(n4160), .Y(n4294) );
  NOR3XLTS U4203 ( .A(rege_out[1]), .B(rege_out[0]), .C(n3961), .Y(n3989) );
  NAND2X1TS U4204 ( .A(n3989), .B(n4812), .Y(n4157) );
  INVX2TS U4205 ( .A(counterii[1]), .Y(n4418) );
  NAND2X1TS U4206 ( .A(ssr_ms0[1]), .B(n4418), .Y(n3265) );
  INVX2TS U4207 ( .A(ssr_ms0[0]), .Y(n3751) );
  OR2X1TS U4208 ( .A(n3265), .B(n3751), .Y(n4126) );
  NOR3BX2TS U4209 ( .AN(mux12[1]), .B(mux12[0]), .C(n3276), .Y(n4293) );
  INVX2TS U4210 ( .A(n3271), .Y(n3273) );
  OAI22X1TS U4211 ( .A0(alu1[1]), .A1(alu1[0]), .B0(n3267), .B1(n3266), .Y(
        n3272) );
  OAI32X1TS U4212 ( .A0(n3268), .A1(n2316), .A2(n3419), .B0(n3355), .B1(n3267), 
        .Y(n3269) );
  OAI32X1TS U4213 ( .A0(n3273), .A1(n3403), .A2(n3272), .B0(n3271), .B1(n3270), 
        .Y(n3274) );
  NOR3XLTS U4214 ( .A(mux12[1]), .B(mux12[0]), .C(n3276), .Y(n3277) );
  BUFX3TS U4215 ( .A(n3277), .Y(n4290) );
  AOI22X1TS U4216 ( .A0(n4293), .A1(aluone_out[0]), .B0(n4290), .B1(
        mult1_out[0]), .Y(n3278) );
  NAND2BXLTS U4217 ( .AN(ssr_ms0[1]), .B(counterii[1]), .Y(n3880) );
  OAI211XLTS U4218 ( .A0(n4300), .A1(n4126), .B0(n3278), .C0(n4135), .Y(n3281)
         );
  INVX2TS U4219 ( .A(count_out[2]), .Y(n3279) );
  INVX2TS U4220 ( .A(count_out[0]), .Y(n3932) );
  INVX2TS U4221 ( .A(count_out[1]), .Y(n3931) );
  AOI31XLTS U4222 ( .A0(n3279), .A1(n3932), .A2(n3931), .B0(n3880), .Y(n4225)
         );
  NOR3XLTS U4223 ( .A(count_out[5]), .B(count_out[4]), .C(n3880), .Y(n4171) );
  INVX2TS U4224 ( .A(count_out[3]), .Y(n4075) );
  OAI21XLTS U4225 ( .A0(ssr_ms0[1]), .A1(ssr_ms0[0]), .B0(n4418), .Y(n3934) );
  INVX2TS U4226 ( .A(n3934), .Y(n4170) );
  AOI21X1TS U4227 ( .A0(n4171), .A1(n4075), .B0(n4170), .Y(n4291) );
  NOR2XLTS U4228 ( .A(n4225), .B(n4291), .Y(n3280) );
  MXI2XLTS U4229 ( .A(ssrms0_out[0]), .B(n3281), .S0(n3280), .Y(n3282) );
  OAI21XLTS U4230 ( .A0(n4294), .A1(n4157), .B0(n3282), .Y(n1879) );
  NAND2X1TS U4231 ( .A(sr_res[0]), .B(sr_res[1]), .Y(n3299) );
  INVX2TS U4232 ( .A(regres_out[2]), .Y(n4642) );
  NOR2XLTS U4233 ( .A(sr_res[0]), .B(n4603), .Y(n4598) );
  INVX2TS U4234 ( .A(n4598), .Y(n3441) );
  INVX2TS U4235 ( .A(n3441), .Y(n3723) );
  AOI22X1TS U4236 ( .A0(regres_out[1]), .A1(n4603), .B0(regres_out[0]), .B1(
        n3723), .Y(n3285) );
  NAND2BXLTS U4237 ( .AN(sr_res[1]), .B(sr_res[0]), .Y(n3346) );
  NOR2XLTS U4238 ( .A(mux21[0]), .B(n3346), .Y(n3345) );
  OAI2BB2XLTS U4239 ( .B0(mux21[1]), .B1(n3346), .A0N(n3345), .A1N(n_input[1]), 
        .Y(n3283) );
  OAI31X1TS U4240 ( .A0(mux21[0]), .A1(mux21[1]), .A2(aluone_out[1]), .B0(
        n3283), .Y(n3284) );
  OAI211XLTS U4241 ( .A0(n3299), .A1(n4642), .B0(n3285), .C0(n3284), .Y(n1688)
         );
  INVX2TS U4242 ( .A(mux14[0]), .Y(n4746) );
  NOR2X1TS U4243 ( .A(n4746), .B(n1991), .Y(n4771) );
  INVX2TS U4244 ( .A(n4771), .Y(n4750) );
  NAND2X1TS U4245 ( .A(n1991), .B(mux14[0]), .Y(n4749) );
  INVX2TS U4246 ( .A(n4749), .Y(n4769) );
  AOI22X1TS U4247 ( .A0(n3286), .A1(srmq_out[32]), .B0(n4769), .B1(
        calculator_input[9]), .Y(n3287) );
  OAI21XLTS U4248 ( .A0(n4750), .A1(n3288), .B0(n3287), .Y(m14_out[9]) );
  AOI22X1TS U4249 ( .A0(n3286), .A1(srmq_out[31]), .B0(n4769), .B1(
        calculator_input[8]), .Y(n3289) );
  OAI21XLTS U4250 ( .A0(n4750), .A1(n3290), .B0(n3289), .Y(m14_out[8]) );
  AOI22X1TS U4251 ( .A0(n3286), .A1(srmq_out[37]), .B0(n4769), .B1(
        calculator_input[14]), .Y(n3291) );
  OAI21XLTS U4252 ( .A0(n4750), .A1(n3292), .B0(n3291), .Y(m14_out[14]) );
  AOI22X1TS U4253 ( .A0(n3286), .A1(srmq_out[39]), .B0(n4769), .B1(
        calculator_input[16]), .Y(n3293) );
  OAI21XLTS U4254 ( .A0(n4750), .A1(n3294), .B0(n3293), .Y(m14_out[16]) );
  AOI22X1TS U4255 ( .A0(n3286), .A1(srmq_out[27]), .B0(n4769), .B1(
        calculator_input[4]), .Y(n3295) );
  OAI21XLTS U4256 ( .A0(n4750), .A1(n3296), .B0(n3295), .Y(m14_out[4]) );
  AOI22X1TS U4257 ( .A0(n3286), .A1(srmq_out[42]), .B0(n4769), .B1(
        calculator_input[19]), .Y(n3297) );
  OAI21XLTS U4258 ( .A0(n4750), .A1(n3298), .B0(n3297), .Y(m14_out[19]) );
  INVX2TS U4259 ( .A(aluone_out[2]), .Y(n4283) );
  NOR3XLTS U4260 ( .A(mux21[0]), .B(mux21[1]), .C(n3346), .Y(n4601) );
  INVX2TS U4261 ( .A(n4601), .Y(n3726) );
  INVX2TS U4262 ( .A(n3299), .Y(n4604) );
  AOI22X1TS U4263 ( .A0(regres_out[3]), .A1(n4604), .B0(regres_out[2]), .B1(
        n4603), .Y(n3301) );
  CLKAND2X2TS U4264 ( .A(n3345), .B(mux21[1]), .Y(n4602) );
  AOI22X1TS U4265 ( .A0(regres_out[1]), .A1(n3723), .B0(n4602), .B1(n_input[2]), .Y(n3300) );
  OAI211XLTS U4266 ( .A0(n4283), .A1(n3726), .B0(n3301), .C0(n3300), .Y(n1689)
         );
  AOI32X1TS U4267 ( .A0(n4715), .A1(n4722), .A2(n3497), .B0(m18_out[0]), .B1(
        n4722), .Y(n3307) );
  NAND2X1TS U4268 ( .A(m18_out[0]), .B(m17_out[0]), .Y(n3302) );
  OAI22X1TS U4269 ( .A0(n3501), .A1(n3303), .B0(n3302), .B1(n3503), .Y(n3304)
         );
  AOI21X1TS U4270 ( .A0(n3307), .A1(m17_out[0]), .B0(n3304), .Y(n3305) );
  OAI31X1TS U4271 ( .A0(n3307), .A1(n3306), .A2(m17_out[0]), .B0(n3305), .Y(
        alutwo_out[0]) );
  INVX2TS U4272 ( .A(n4741), .Y(n3343) );
  AOI22X1TS U4273 ( .A0(n4740), .A1(alutwo_out[0]), .B0(n3343), .B1(
        rf_aout[23]), .Y(n3308) );
  NAND2X1TS U4274 ( .A(mux13[0]), .B(n3343), .Y(n3389) );
  OAI211XLTS U4275 ( .A0(n3159), .A1(n4785), .B0(n3308), .C0(n3389), .Y(
        m3_out[23]) );
  INVX2TS U4276 ( .A(n3309), .Y(n3313) );
  NAND2X1TS U4277 ( .A(n4689), .B(n3320), .Y(n3314) );
  AOI32X1TS U4278 ( .A0(n3503), .A1(m18_out[2]), .A2(n3314), .B0(n3311), .B1(
        n3310), .Y(n3312) );
  AOI21X1TS U4279 ( .A0(n3445), .A1(n4710), .B0(n2455), .Y(n3342) );
  OAI32X1TS U4280 ( .A0(m17_out[2]), .A1(m18_out[2]), .A2(n3314), .B0(n3342), 
        .B1(m17_out[2]), .Y(n3315) );
  AOI21X1TS U4281 ( .A0(n3316), .A1(n3493), .B0(n3315), .Y(n3324) );
  NOR2BX1TS U4282 ( .AN(n3318), .B(n3317), .Y(n3319) );
  XNOR2X1TS U4283 ( .A(m18_out[2]), .B(n3319), .Y(n3322) );
  OAI31X1TS U4284 ( .A0(m17_out[2]), .A1(n4715), .A2(n3320), .B0(n3501), .Y(
        n3321) );
  AOI22X1TS U4285 ( .A0(n3322), .A1(n3499), .B0(m18_out[2]), .B1(n3321), .Y(
        n3323) );
  AOI22X1TS U4286 ( .A0(n4740), .A1(alutwo_out[2]), .B0(n3343), .B1(
        rf_aout[25]), .Y(n3327) );
  OAI211XLTS U4287 ( .A0(n3159), .A1(n4781), .B0(n3327), .C0(n3389), .Y(
        m3_out[25]) );
  AOI22X1TS U4288 ( .A0(n4740), .A1(alutwo_out[1]), .B0(n3343), .B1(
        rf_aout[24]), .Y(n3328) );
  OAI211XLTS U4289 ( .A0(n3159), .A1(n4775), .B0(n3328), .C0(n3389), .Y(
        m3_out[24]) );
  AOI22X1TS U4290 ( .A0(n3493), .A1(n3330), .B0(m17_out[3]), .B1(n3329), .Y(
        n3341) );
  NOR2BX1TS U4291 ( .AN(n3332), .B(n3331), .Y(n3334) );
  OAI22X1TS U4292 ( .A0(n3334), .A1(n3497), .B0(n4715), .B1(n3335), .Y(n3338)
         );
  AOI22X1TS U4293 ( .A0(n4689), .A1(n3335), .B0(n3499), .B1(n3334), .Y(n3336)
         );
  AOI22X1TS U4294 ( .A0(n3339), .A1(n3338), .B0(n3337), .B1(m18_out[3]), .Y(
        n3340) );
  AOI22X1TS U4295 ( .A0(n4740), .A1(alutwo_out[3]), .B0(n3343), .B1(
        rf_aout[26]), .Y(n3344) );
  OAI211XLTS U4296 ( .A0(n3159), .A1(n4782), .B0(n3344), .C0(n3389), .Y(
        m3_out[26]) );
  AOI22X1TS U4297 ( .A0(regres_out[4]), .A1(n4604), .B0(regres_out[3]), .B1(
        n4603), .Y(n3349) );
  OAI2BB2XLTS U4298 ( .B0(mux21[1]), .B1(n3346), .A0N(n3345), .A1N(n_input[3]), 
        .Y(n3347) );
  OAI31X1TS U4299 ( .A0(mux21[0]), .A1(mux21[1]), .A2(aluone_out[3]), .B0(
        n3347), .Y(n3348) );
  OAI211XLTS U4300 ( .A0(n3441), .A1(n4642), .B0(n3349), .C0(n3348), .Y(n1690)
         );
  AOI22X1TS U4301 ( .A0(n3361), .A1(n3403), .B0(n3360), .B1(n3359), .Y(n3368)
         );
  OAI22X1TS U4302 ( .A0(n3363), .A1(n3739), .B0(n3741), .B1(n3362), .Y(n3364)
         );
  AOI22X1TS U4303 ( .A0(n3366), .A1(n3365), .B0(n3370), .B1(n3364), .Y(n3367)
         );
  INVX2TS U4304 ( .A(aluone_out[4]), .Y(n4262) );
  AOI22X1TS U4305 ( .A0(regres_out[5]), .A1(n4604), .B0(regres_out[4]), .B1(
        n4603), .Y(n3372) );
  AOI22X1TS U4306 ( .A0(regres_out[3]), .A1(n3723), .B0(n4602), .B1(n_input[4]), .Y(n3371) );
  OAI211XLTS U4307 ( .A0(n4262), .A1(n3726), .B0(n3372), .C0(n3371), .Y(n1691)
         );
  INVX2TS U4308 ( .A(rf_aout[28]), .Y(n3481) );
  NOR2BX1TS U4309 ( .AN(n3376), .B(n3375), .Y(n3380) );
  OA22X1TS U4310 ( .A0(n4715), .A1(n3381), .B0(n3497), .B1(n3380), .Y(n3388)
         );
  INVX2TS U4311 ( .A(m17_out[5]), .Y(n3383) );
  AOI21X1TS U4312 ( .A0(n4710), .A1(n3378), .B0(n3526), .Y(n3379) );
  AOI22X1TS U4313 ( .A0(n4689), .A1(n3381), .B0(n3499), .B1(n3380), .Y(n3382)
         );
  AOI22X1TS U4314 ( .A0(n3493), .A1(n3385), .B0(m18_out[5]), .B1(n3384), .Y(
        n3386) );
  AOI22X1TS U4315 ( .A0(n4740), .A1(alutwo_out[5]), .B0(n4739), .B1(
        regsum_out[28]), .Y(n3390) );
  OAI211XLTS U4316 ( .A0(n4741), .A1(n3481), .B0(n3390), .C0(n3389), .Y(
        m3_out[28]) );
  INVX2TS U4317 ( .A(aluone_out[5]), .Y(n4253) );
  AOI22X1TS U4318 ( .A0(regres_out[6]), .A1(n4604), .B0(regres_out[5]), .B1(
        n4603), .Y(n3392) );
  AOI22X1TS U4319 ( .A0(regres_out[4]), .A1(n3723), .B0(n4602), .B1(n_input[5]), .Y(n3391) );
  OAI211XLTS U4320 ( .A0(n4253), .A1(n3726), .B0(n3392), .C0(n3391), .Y(n1692)
         );
  INVX2TS U4321 ( .A(aluone_out[6]), .Y(n4244) );
  AOI22X1TS U4322 ( .A0(regres_out[7]), .A1(n4604), .B0(regres_out[6]), .B1(
        n4603), .Y(n3394) );
  AOI22X1TS U4323 ( .A0(regres_out[5]), .A1(n3723), .B0(n4602), .B1(n_input[6]), .Y(n3393) );
  OAI211XLTS U4324 ( .A0(n4244), .A1(n3726), .B0(n3394), .C0(n3393), .Y(n1693)
         );
  OAI2BB2XLTS U4325 ( .B0(n3426), .B1(n3396), .A0N(n3396), .A1N(n3426), .Y(
        n3399) );
  AOI22X1TS U4326 ( .A0(n3398), .A1(n3397), .B0(n3425), .B1(n3426), .Y(n3406)
         );
  AOI22X1TS U4327 ( .A0(n3419), .A1(n3399), .B0(n3736), .B1(n3426), .Y(n3400)
         );
  AOI22X1TS U4328 ( .A0(n3404), .A1(n3403), .B0(n3407), .B1(n3402), .Y(n3405)
         );
  INVX2TS U4329 ( .A(aluone_out[7]), .Y(n4236) );
  AOI22X1TS U4330 ( .A0(regres_out[8]), .A1(n4604), .B0(regres_out[7]), .B1(
        n4603), .Y(n3410) );
  AOI22X1TS U4331 ( .A0(regres_out[6]), .A1(n3723), .B0(n4602), .B1(n_input[7]), .Y(n3409) );
  OAI211XLTS U4332 ( .A0(n4236), .A1(n3726), .B0(n3410), .C0(n3409), .Y(n1694)
         );
  AOI22X1TS U4333 ( .A0(n3411), .A1(rf_aout[30]), .B0(n4740), .B1(
        alutwo_out[7]), .Y(n3412) );
  OAI21XLTS U4334 ( .A0(n3159), .A1(n4783), .B0(n3412), .Y(m3_out[30]) );
  AOI222XLTS U4335 ( .A0(n1991), .A1(n4746), .B0(n1991), .B1(
        calculator_input[23]), .C0(n4746), .C1(alutwo_out[0]), .Y(n3413) );
  OAI21XLTS U4336 ( .A0(n4750), .A1(n3414), .B0(n3413), .Y(m14_out[23]) );
  AOI222XLTS U4337 ( .A0(n1991), .A1(n4746), .B0(n1991), .B1(
        calculator_input[25]), .C0(n4746), .C1(alutwo_out[2]), .Y(n3415) );
  OAI21XLTS U4338 ( .A0(n4750), .A1(n3416), .B0(n3415), .Y(m14_out[25]) );
  AOI22X1TS U4339 ( .A0(regres_out[9]), .A1(n4604), .B0(regres_out[8]), .B1(
        n4603), .Y(n3440) );
  NOR2BX1TS U4340 ( .AN(n3418), .B(n3417), .Y(n3421) );
  AOI21X1TS U4341 ( .A0(n3421), .A1(n3427), .B0(n3420), .Y(n3438) );
  AOI21X1TS U4342 ( .A0(n3729), .A1(n3426), .B0(n3425), .Y(n3430) );
  OAI22X1TS U4343 ( .A0(n3431), .A1(n3430), .B0(n3429), .B1(n3739), .Y(n3436)
         );
  OAI22X1TS U4344 ( .A0(n3434), .A1(n3433), .B0(n3748), .B1(n3432), .Y(n3435)
         );
  OR4X2TS U4345 ( .A(n3438), .B(n3437), .C(n3436), .D(n3435), .Y(aluone_out[8]) );
  AOI22X1TS U4346 ( .A0(n4602), .A1(n_input[8]), .B0(n4601), .B1(aluone_out[8]), .Y(n3439) );
  OAI211XLTS U4347 ( .A0(n3442), .A1(n3441), .B0(n3440), .C0(n3439), .Y(n1695)
         );
  AOI222XLTS U4348 ( .A0(n1991), .A1(n4746), .B0(n1991), .B1(
        calculator_input[26]), .C0(n4746), .C1(alutwo_out[3]), .Y(n3443) );
  OAI21XLTS U4349 ( .A0(n4750), .A1(n3444), .B0(n3443), .Y(m14_out[26]) );
  AOI32X1TS U4350 ( .A0(n3446), .A1(n4722), .A2(n3445), .B0(n4660), .B1(n4722), 
        .Y(n3447) );
  AOI22X1TS U4351 ( .A0(n3493), .A1(n3448), .B0(m17_out[4]), .B1(n3447), .Y(
        n3461) );
  NOR2BX1TS U4352 ( .AN(n3450), .B(n3449), .Y(n3453) );
  OAI22X1TS U4353 ( .A0(n3453), .A1(n3497), .B0(n4715), .B1(n3454), .Y(n3458)
         );
  AOI22X1TS U4354 ( .A0(n4689), .A1(n3454), .B0(n3499), .B1(n3453), .Y(n3455)
         );
  AOI22X1TS U4355 ( .A0(n3459), .A1(n3458), .B0(n3457), .B1(m18_out[4]), .Y(
        n3460) );
  INVX2TS U4356 ( .A(aluone_out[9]), .Y(n3465) );
  AOI22X1TS U4357 ( .A0(regres_out[10]), .A1(n4604), .B0(regres_out[9]), .B1(
        n4603), .Y(n3464) );
  AOI22X1TS U4358 ( .A0(regres_out[8]), .A1(n3723), .B0(n4602), .B1(n_input[9]), .Y(n3463) );
  OAI211XLTS U4359 ( .A0(n3465), .A1(n3726), .B0(n3464), .C0(n3463), .Y(n1696)
         );
  INVX2TS U4360 ( .A(aluone_out[10]), .Y(n4210) );
  AOI22X1TS U4361 ( .A0(regres_out[11]), .A1(n4604), .B0(regres_out[10]), .B1(
        n4603), .Y(n3467) );
  AOI22X1TS U4362 ( .A0(regres_out[9]), .A1(n3723), .B0(n4602), .B1(
        n_input[10]), .Y(n3466) );
  OAI211XLTS U4363 ( .A0(n4210), .A1(n3726), .B0(n3467), .C0(n3466), .Y(n1697)
         );
  INVX2TS U4364 ( .A(aluone_out[11]), .Y(n4201) );
  AOI22X1TS U4365 ( .A0(regres_out[12]), .A1(n4604), .B0(regres_out[11]), .B1(
        n4603), .Y(n3469) );
  AOI22X1TS U4366 ( .A0(regres_out[10]), .A1(n3723), .B0(n4602), .B1(
        n_input[11]), .Y(n3468) );
  OAI211XLTS U4367 ( .A0(n4201), .A1(n3726), .B0(n3469), .C0(n3468), .Y(n1698)
         );
  AOI21X1TS U4368 ( .A0(n3471), .A1(n3470), .B0(n4713), .Y(n3479) );
  INVX2TS U4369 ( .A(n4718), .Y(n3478) );
  NAND2X1TS U4370 ( .A(n4717), .B(n4714), .Y(n3473) );
  OAI22X1TS U4371 ( .A0(n3476), .A1(n3475), .B0(n3474), .B1(n3473), .Y(n3477)
         );
  AOI222XLTS U4372 ( .A0(n1991), .A1(n4746), .B0(n1991), .B1(
        calculator_input[28]), .C0(n4746), .C1(alutwo_out[5]), .Y(n3480) );
  OAI21XLTS U4373 ( .A0(n4750), .A1(n3481), .B0(n3480), .Y(m14_out[28]) );
  OAI2BB2XLTS U4374 ( .B0(n3482), .B1(n4660), .A0N(n4689), .A1N(n3483), .Y(
        n3485) );
  OAI32X1TS U4375 ( .A0(n3486), .A1(n3526), .A2(n3485), .B0(m17_out[10]), .B1(
        n3484), .Y(n3489) );
  AOI32X1TS U4376 ( .A0(n3487), .A1(n4696), .A2(n4711), .B0(n3518), .B1(n4696), 
        .Y(n3488) );
  AOI22X1TS U4377 ( .A0(n3493), .A1(n3492), .B0(m17_out[6]), .B1(n3491), .Y(
        n3509) );
  NOR2BX1TS U4378 ( .AN(n3495), .B(n3494), .Y(n3498) );
  OAI22X1TS U4379 ( .A0(n3498), .A1(n3497), .B0(n4715), .B1(n3500), .Y(n3506)
         );
  AOI22X1TS U4380 ( .A0(n4689), .A1(n3500), .B0(n3499), .B1(n3498), .Y(n3502)
         );
  AOI22X1TS U4381 ( .A0(n3507), .A1(n3506), .B0(n3505), .B1(m18_out[6]), .Y(
        n3508) );
  AOI222XLTS U4382 ( .A0(n1991), .A1(n4746), .B0(n1991), .B1(
        calculator_input[29]), .C0(n4746), .C1(alutwo_out[6]), .Y(n3511) );
  OAI21XLTS U4383 ( .A0(n4750), .A1(n4737), .B0(n3511), .Y(m14_out[29]) );
  AOI22X1TS U4384 ( .A0(calculator_input[30]), .A1(n4769), .B0(n3286), .B1(
        alutwo_out[7]), .Y(n3512) );
  OAI21XLTS U4385 ( .A0(n3513), .A1(n4750), .B0(n3512), .Y(m14_out[30]) );
  INVX2TS U4386 ( .A(aluone_out[12]), .Y(n3516) );
  AOI22X1TS U4387 ( .A0(regres_out[13]), .A1(n4604), .B0(regres_out[12]), .B1(
        n4603), .Y(n3515) );
  AOI22X1TS U4388 ( .A0(regres_out[11]), .A1(n3723), .B0(n4602), .B1(
        n_input[12]), .Y(n3514) );
  OAI211XLTS U4389 ( .A0(n3516), .A1(n3726), .B0(n3515), .C0(n3514), .Y(n1699)
         );
  OA21XLTS U4390 ( .A0(n3518), .A1(n3517), .B0(n3530), .Y(n3525) );
  OAI2BB2XLTS U4391 ( .B0(n3548), .B1(n4715), .A0N(n4710), .A1N(n3520), .Y(
        n3522) );
  NAND2X1TS U4392 ( .A(n4689), .B(n3548), .Y(n3519) );
  OAI32X1TS U4393 ( .A0(n3523), .A1(n3526), .A2(n3522), .B0(m17_out[11]), .B1(
        n3521), .Y(n3524) );
  AOI21X1TS U4394 ( .A0(n4689), .A1(n3527), .B0(n3526), .Y(n3549) );
  AOI21X1TS U4395 ( .A0(m17_out[12]), .A1(n3529), .B0(n4700), .Y(n3533) );
  AOI32X1TS U4396 ( .A0(n3531), .A1(n4696), .A2(n3530), .B0(n4699), .B1(n4696), 
        .Y(n3532) );
  INVX2TS U4397 ( .A(aluone_out[13]), .Y(n3537) );
  AOI22X1TS U4398 ( .A0(regres_out[14]), .A1(n4604), .B0(regres_out[13]), .B1(
        n4603), .Y(n3536) );
  AOI22X1TS U4399 ( .A0(regres_out[12]), .A1(n3723), .B0(n4602), .B1(
        n_input[13]), .Y(n3535) );
  OAI211XLTS U4400 ( .A0(n3537), .A1(n3726), .B0(n3536), .C0(n3535), .Y(n1700)
         );
  AOI21X1TS U4401 ( .A0(n3538), .A1(n3545), .B0(n4685), .Y(n3544) );
  OA21XLTS U4402 ( .A0(n3539), .A1(n4660), .B0(n4722), .Y(n4693) );
  OAI32X1TS U4403 ( .A0(m17_out[16]), .A1(n2455), .A2(n3542), .B0(n3541), .B1(
        n3540), .Y(n3543) );
  OA21XLTS U4404 ( .A0(n3561), .A1(n3546), .B0(n3545), .Y(n3555) );
  OAI22X1TS U4405 ( .A0(n3550), .A1(n4701), .B0(n4660), .B1(n3565), .Y(n3553)
         );
  INVX2TS U4406 ( .A(n3549), .Y(n4702) );
  AOI21X1TS U4407 ( .A0(n4689), .A1(n3550), .B0(n4702), .Y(n3556) );
  OAI2BB1X1TS U4408 ( .A0N(n3565), .A1N(n4710), .B0(n3556), .Y(n3551) );
  OAI32X1TS U4409 ( .A0(m17_out[15]), .A1(n2455), .A2(n3553), .B0(n3552), .B1(
        n3551), .Y(n3554) );
  AOI22X1TS U4410 ( .A0(n3560), .A1(n3559), .B0(n3558), .B1(m17_out[14]), .Y(
        n3564) );
  AOI32X1TS U4411 ( .A0(n3562), .A1(n4696), .A2(n4697), .B0(n3561), .B1(n4696), 
        .Y(n3563) );
  INVX2TS U4412 ( .A(aluone_out[14]), .Y(n3568) );
  AOI22X1TS U4413 ( .A0(regres_out[15]), .A1(n4604), .B0(regres_out[14]), .B1(
        n4603), .Y(n3567) );
  AOI22X1TS U4414 ( .A0(regres_out[13]), .A1(n3723), .B0(n4602), .B1(
        n_input[14]), .Y(n3566) );
  OAI211XLTS U4415 ( .A0(n3568), .A1(n3726), .B0(n3567), .C0(n3566), .Y(n1701)
         );
  AOI21X1TS U4416 ( .A0(n3570), .A1(n4683), .B0(n3569), .Y(n3577) );
  NAND2X1TS U4417 ( .A(n4710), .B(n3571), .Y(n3572) );
  OAI32X1TS U4418 ( .A0(m17_out[18]), .A1(n3575), .A2(n4687), .B0(n3574), .B1(
        n3573), .Y(n3576) );
  INVX2TS U4419 ( .A(aluone_out[15]), .Y(n3580) );
  AOI22X1TS U4420 ( .A0(regres_out[16]), .A1(n4604), .B0(regres_out[15]), .B1(
        n4603), .Y(n3579) );
  AOI22X1TS U4421 ( .A0(regres_out[14]), .A1(n3723), .B0(n4602), .B1(
        n_input[15]), .Y(n3578) );
  OAI211XLTS U4422 ( .A0(n3580), .A1(n3726), .B0(n3579), .C0(n3578), .Y(n1702)
         );
  INVX2TS U4423 ( .A(aluone_out[16]), .Y(n4161) );
  AOI22X1TS U4424 ( .A0(regres_out[17]), .A1(n4604), .B0(regres_out[16]), .B1(
        n4603), .Y(n3582) );
  AOI22X1TS U4425 ( .A0(regres_out[15]), .A1(n3723), .B0(n4602), .B1(
        n_input[16]), .Y(n3581) );
  OAI211XLTS U4426 ( .A0(n4161), .A1(n3726), .B0(n3582), .C0(n3581), .Y(n1703)
         );
  AOI21X1TS U4427 ( .A0(n3584), .A1(n3583), .B0(n3597), .Y(n3592) );
  AOI32X1TS U4428 ( .A0(n4710), .A1(n3590), .A2(n3589), .B0(n3588), .B1(n3590), 
        .Y(n3591) );
  AOI21X1TS U4429 ( .A0(n4689), .A1(n3595), .B0(n3594), .Y(n3610) );
  AOI22X1TS U4430 ( .A0(n3611), .A1(n3599), .B0(n4696), .B1(n3598), .Y(n3601)
         );
  INVX2TS U4431 ( .A(aluone_out[17]), .Y(n3604) );
  AOI22X1TS U4432 ( .A0(regres_out[18]), .A1(n4604), .B0(regres_out[17]), .B1(
        n4603), .Y(n3603) );
  AOI22X1TS U4433 ( .A0(regres_out[16]), .A1(n3723), .B0(n4602), .B1(
        n_input[17]), .Y(n3602) );
  OAI211XLTS U4434 ( .A0(n3604), .A1(n3726), .B0(n3603), .C0(n3602), .Y(n1704)
         );
  AOI21X1TS U4435 ( .A0(n3606), .A1(n3605), .B0(n3621), .Y(n3614) );
  INVX2TS U4436 ( .A(aluone_out[18]), .Y(n4129) );
  AOI22X1TS U4437 ( .A0(regres_out[19]), .A1(n4604), .B0(regres_out[18]), .B1(
        n4603), .Y(n3616) );
  AOI22X1TS U4438 ( .A0(regres_out[17]), .A1(n3723), .B0(n4602), .B1(
        n_input[18]), .Y(n3615) );
  OAI211XLTS U4439 ( .A0(n4129), .A1(n3726), .B0(n3616), .C0(n3615), .Y(n1705)
         );
  OAI31X1TS U4440 ( .A0(n3619), .A1(n2455), .A2(n3618), .B0(n3617), .Y(n3625)
         );
  INVX2TS U4441 ( .A(n3634), .Y(n4678) );
  AOI22X1TS U4442 ( .A0(n4696), .A1(n3623), .B0(m17_out[23]), .B1(n4678), .Y(
        n3624) );
  OA21XLTS U4443 ( .A0(n4670), .A1(n3626), .B0(n3636), .Y(n3633) );
  OAI22X1TS U4444 ( .A0(n3627), .A1(n4660), .B0(n4715), .B1(m17_out[24]), .Y(
        n3629) );
  NAND2X1TS U4445 ( .A(n4689), .B(n3645), .Y(n4673) );
  OAI32X1TS U4446 ( .A0(n3630), .A1(n4678), .A2(n3629), .B0(n3628), .B1(
        m17_out[25]), .Y(n3632) );
  INVX2TS U4447 ( .A(n3639), .Y(n4677) );
  INVX2TS U4448 ( .A(n3638), .Y(n3635) );
  NAND2X1TS U4449 ( .A(n4677), .B(n3635), .Y(n3631) );
  AOI21X1TS U4450 ( .A0(n4689), .A1(n3665), .B0(n3669), .Y(n3648) );
  AOI32X1TS U4451 ( .A0(n3637), .A1(n4696), .A2(n3636), .B0(n3647), .B1(n4696), 
        .Y(n3643) );
  NAND2X1TS U4452 ( .A(m17_out[24]), .B(m17_out[25]), .Y(n3640) );
  OAI22X1TS U4453 ( .A0(n3640), .A1(n4673), .B0(n3639), .B1(n3638), .Y(n3641)
         );
  INVX2TS U4454 ( .A(n3665), .Y(n3644) );
  AOI22X1TS U4455 ( .A0(n4696), .A1(n3651), .B0(m17_out[27]), .B1(n3650), .Y(
        n3653) );
  NAND2X1TS U4456 ( .A(n4677), .B(n3671), .Y(n3652) );
  INVX2TS U4457 ( .A(aluone_out[20]), .Y(n3657) );
  AOI22X1TS U4458 ( .A0(regres_out[21]), .A1(n4604), .B0(regres_out[20]), .B1(
        n4603), .Y(n3656) );
  AOI22X1TS U4459 ( .A0(regres_out[19]), .A1(n3723), .B0(n4602), .B1(
        n_input[20]), .Y(n3655) );
  OAI211XLTS U4460 ( .A0(n3657), .A1(n3726), .B0(n3656), .C0(n3655), .Y(n1707)
         );
  INVX2TS U4461 ( .A(aluone_out[19]), .Y(n3660) );
  AOI22X1TS U4462 ( .A0(regres_out[20]), .A1(n4604), .B0(regres_out[19]), .B1(
        n4603), .Y(n3659) );
  AOI22X1TS U4463 ( .A0(regres_out[18]), .A1(n3723), .B0(n4602), .B1(
        n_input[19]), .Y(n3658) );
  OAI211XLTS U4464 ( .A0(n3660), .A1(n3726), .B0(n3659), .C0(n3658), .Y(n1706)
         );
  AOI21X1TS U4465 ( .A0(n3662), .A1(n3661), .B0(n3678), .Y(n3673) );
  OAI22X1TS U4466 ( .A0(n3664), .A1(n4715), .B0(n3663), .B1(n4660), .Y(n3668)
         );
  OAI31X1TS U4467 ( .A0(n3666), .A1(n3665), .A2(n4673), .B0(n4714), .Y(n3667)
         );
  OAI32X1TS U4468 ( .A0(n3670), .A1(n3669), .A2(n3668), .B0(n3667), .B1(
        m17_out[28]), .Y(n3672) );
  INVX2TS U4469 ( .A(aluone_out[21]), .Y(n4093) );
  AOI22X1TS U4470 ( .A0(regres_out[22]), .A1(n4604), .B0(regres_out[21]), .B1(
        n4603), .Y(n3675) );
  AOI22X1TS U4471 ( .A0(regres_out[20]), .A1(n3723), .B0(n4602), .B1(
        n_input[21]), .Y(n3674) );
  OAI211XLTS U4472 ( .A0(n4093), .A1(n3726), .B0(n3675), .C0(n3674), .Y(n1708)
         );
  OA21XLTS U4473 ( .A0(n3678), .A1(n3677), .B0(n3676), .Y(n3689) );
  INVX2TS U4474 ( .A(n3679), .Y(n3681) );
  OAI31X1TS U4475 ( .A0(n2455), .A1(n3682), .A2(n3681), .B0(n3680), .Y(n3688)
         );
  AOI21X1TS U4476 ( .A0(n4689), .A1(n3684), .B0(n3683), .Y(n3696) );
  INVX2TS U4477 ( .A(n3696), .Y(n3685) );
  AOI32X1TS U4478 ( .A0(n4710), .A1(m17_out[29]), .A2(n3686), .B0(n3685), .B1(
        m17_out[29]), .Y(n3687) );
  XNOR2X1TS U4479 ( .A(n3692), .B(n3691), .Y(n3701) );
  OAI31X1TS U4480 ( .A0(n3695), .A1(n3694), .A2(n2455), .B0(n3693), .Y(n3700)
         );
  OAI2BB2XLTS U4481 ( .B0(m17_out[30]), .B1(n4715), .A0N(n4710), .A1N(n3697), 
        .Y(n3698) );
  INVX2TS U4482 ( .A(aluone_out[22]), .Y(n3704) );
  AOI22X1TS U4483 ( .A0(regres_out[23]), .A1(n4604), .B0(regres_out[22]), .B1(
        n4603), .Y(n3703) );
  AOI22X1TS U4484 ( .A0(regres_out[21]), .A1(n3723), .B0(n4602), .B1(
        n_input[22]), .Y(n3702) );
  OAI211XLTS U4485 ( .A0(n3704), .A1(n3726), .B0(n3703), .C0(n3702), .Y(n1709)
         );
  INVX2TS U4486 ( .A(aluone_out[23]), .Y(n4071) );
  AOI22X1TS U4487 ( .A0(regres_out[24]), .A1(n4604), .B0(regres_out[23]), .B1(
        n4603), .Y(n3706) );
  AOI22X1TS U4488 ( .A0(regres_out[22]), .A1(n3723), .B0(n4602), .B1(
        n_input[23]), .Y(n3705) );
  OAI211XLTS U4489 ( .A0(n4071), .A1(n3726), .B0(n3706), .C0(n3705), .Y(n1710)
         );
  INVX2TS U4490 ( .A(aluone_out[24]), .Y(n4059) );
  AOI22X1TS U4491 ( .A0(regres_out[25]), .A1(n4604), .B0(regres_out[24]), .B1(
        n4603), .Y(n3708) );
  AOI22X1TS U4492 ( .A0(regres_out[23]), .A1(n3723), .B0(n4602), .B1(
        n_input[24]), .Y(n3707) );
  OAI211XLTS U4493 ( .A0(n4059), .A1(n3726), .B0(n3708), .C0(n3707), .Y(n1711)
         );
  INVX2TS U4494 ( .A(aluone_out[26]), .Y(n3711) );
  AOI22X1TS U4495 ( .A0(regres_out[27]), .A1(n4604), .B0(regres_out[26]), .B1(
        n4603), .Y(n3710) );
  AOI22X1TS U4496 ( .A0(regres_out[25]), .A1(n3723), .B0(n4602), .B1(
        n_input[26]), .Y(n3709) );
  OAI211XLTS U4497 ( .A0(n3711), .A1(n3726), .B0(n3710), .C0(n3709), .Y(n1713)
         );
  INVX2TS U4498 ( .A(aluone_out[25]), .Y(n3714) );
  AOI22X1TS U4499 ( .A0(regres_out[26]), .A1(n4604), .B0(regres_out[25]), .B1(
        n4603), .Y(n3713) );
  AOI22X1TS U4500 ( .A0(regres_out[24]), .A1(n3723), .B0(n4602), .B1(
        n_input[25]), .Y(n3712) );
  OAI211XLTS U4501 ( .A0(n3714), .A1(n3726), .B0(n3713), .C0(n3712), .Y(n1712)
         );
  INVX2TS U4502 ( .A(aluone_out[27]), .Y(n3717) );
  AOI22X1TS U4503 ( .A0(regres_out[28]), .A1(n4604), .B0(regres_out[27]), .B1(
        n4603), .Y(n3716) );
  AOI22X1TS U4504 ( .A0(regres_out[26]), .A1(n3723), .B0(n4602), .B1(
        n_input[27]), .Y(n3715) );
  OAI211XLTS U4505 ( .A0(n3717), .A1(n3726), .B0(n3716), .C0(n3715), .Y(n1714)
         );
  INVX2TS U4506 ( .A(aluone_out[28]), .Y(n4001) );
  AOI22X1TS U4507 ( .A0(regres_out[29]), .A1(n4604), .B0(regres_out[28]), .B1(
        n4603), .Y(n3719) );
  AOI22X1TS U4508 ( .A0(regres_out[27]), .A1(n4598), .B0(n4602), .B1(
        n_input[28]), .Y(n3718) );
  OAI211XLTS U4509 ( .A0(n4001), .A1(n3726), .B0(n3719), .C0(n3718), .Y(n1715)
         );
  INVX2TS U4510 ( .A(aluone_out[30]), .Y(n3722) );
  AOI22X1TS U4511 ( .A0(regres_out[31]), .A1(n4604), .B0(regres_out[30]), .B1(
        n4603), .Y(n3721) );
  AOI22X1TS U4512 ( .A0(regres_out[29]), .A1(n3723), .B0(n4602), .B1(
        n_input[30]), .Y(n3720) );
  OAI211XLTS U4513 ( .A0(n3722), .A1(n3726), .B0(n3721), .C0(n3720), .Y(n1717)
         );
  INVX2TS U4514 ( .A(aluone_out[29]), .Y(n3727) );
  AOI22X1TS U4515 ( .A0(regres_out[30]), .A1(n4604), .B0(regres_out[29]), .B1(
        n4603), .Y(n3725) );
  AOI22X1TS U4516 ( .A0(regres_out[28]), .A1(n3723), .B0(n4602), .B1(
        n_input[29]), .Y(n3724) );
  OAI211XLTS U4517 ( .A0(n3727), .A1(n3726), .B0(n3725), .C0(n3724), .Y(n1716)
         );
  AOI31XLTS U4518 ( .A0(count_out[2]), .A1(count_out[0]), .A2(count_out[1]), 
        .B0(n3880), .Y(n4234) );
  INVX2TS U4519 ( .A(count_out[4]), .Y(n3813) );
  NOR3XLTS U4520 ( .A(count_out[5]), .B(n3880), .C(n3813), .Y(n4076) );
  AOI21X1TS U4521 ( .A0(count_out[3]), .A1(n4076), .B0(n4170), .Y(n4050) );
  NOR2XLTS U4522 ( .A(n4234), .B(n4050), .Y(n3756) );
  INVX2TS U4523 ( .A(ssrms0_out[31]), .Y(n3959) );
  NAND2X1TS U4524 ( .A(n4145), .B(n4778), .Y(n4209) );
  AOI22X1TS U4525 ( .A0(rege_out[0]), .A1(ssrms0_out[16]), .B0(ssrms0_out[17]), 
        .B1(n4811), .Y(n3970) );
  AOI22X1TS U4526 ( .A0(rege_out[0]), .A1(ssrms0_out[18]), .B0(ssrms0_out[19]), 
        .B1(n4811), .Y(n3973) );
  AOI22X1TS U4527 ( .A0(rege_out[1]), .A1(n3970), .B0(n3973), .B1(n4810), .Y(
        n4009) );
  AOI22X1TS U4528 ( .A0(rege_out[0]), .A1(ssrms0_out[20]), .B0(ssrms0_out[21]), 
        .B1(n4811), .Y(n3972) );
  AOI22X1TS U4529 ( .A0(rege_out[0]), .A1(ssrms0_out[22]), .B0(ssrms0_out[23]), 
        .B1(n4811), .Y(n4040) );
  AOI22X1TS U4530 ( .A0(rege_out[1]), .A1(n3972), .B0(n4040), .B1(n4810), .Y(
        n4011) );
  AOI22X1TS U4531 ( .A0(rege_out[2]), .A1(n4009), .B0(n4011), .B1(n4812), .Y(
        n4070) );
  XNOR2X1TS U4532 ( .A(n3733), .B(n3749), .Y(n3740) );
  XNOR2X1TS U4533 ( .A(n3734), .B(n3735), .Y(n3742) );
  AOI22X1TS U4534 ( .A0(n3419), .A1(n3742), .B0(n3736), .B1(n3735), .Y(n3738)
         );
  OAI2BB2XLTS U4535 ( .B0(n3742), .B1(n3741), .A0N(n3740), .A1N(n2316), .Y(
        n3744) );
  INVX2TS U4536 ( .A(n4145), .Y(n4162) );
  NOR2X1TS U4537 ( .A(n4778), .B(n4162), .Y(n4044) );
  AOI22X1TS U4538 ( .A0(rege_out[0]), .A1(ssrms0_out[0]), .B0(ssrms0_out[1]), 
        .B1(n4811), .Y(n3975) );
  AOI22X1TS U4539 ( .A0(rege_out[0]), .A1(ssrms0_out[2]), .B0(ssrms0_out[3]), 
        .B1(n4811), .Y(n3977) );
  AOI22X1TS U4540 ( .A0(rege_out[1]), .A1(n3975), .B0(n3977), .B1(n4810), .Y(
        n4012) );
  AOI22X1TS U4541 ( .A0(rege_out[0]), .A1(ssrms0_out[4]), .B0(ssrms0_out[5]), 
        .B1(n4811), .Y(n3976) );
  AOI22X1TS U4542 ( .A0(rege_out[0]), .A1(ssrms0_out[6]), .B0(ssrms0_out[7]), 
        .B1(n4811), .Y(n3979) );
  AOI22X1TS U4543 ( .A0(rege_out[1]), .A1(n3976), .B0(n3979), .B1(n4810), .Y(
        n4110) );
  AOI22X1TS U4544 ( .A0(rege_out[2]), .A1(n4012), .B0(n4110), .B1(n4812), .Y(
        n4235) );
  AOI22X1TS U4545 ( .A0(rege_out[0]), .A1(ssrms0_out[8]), .B0(ssrms0_out[9]), 
        .B1(n4811), .Y(n3978) );
  AOI22X1TS U4546 ( .A0(rege_out[0]), .A1(ssrms0_out[10]), .B0(ssrms0_out[11]), 
        .B1(n4811), .Y(n3981) );
  AOI22X1TS U4547 ( .A0(rege_out[1]), .A1(n3978), .B0(n3981), .B1(n4810), .Y(
        n4111) );
  AOI22X1TS U4548 ( .A0(rege_out[0]), .A1(ssrms0_out[12]), .B0(ssrms0_out[13]), 
        .B1(n4811), .Y(n3980) );
  AOI22X1TS U4549 ( .A0(rege_out[0]), .A1(ssrms0_out[14]), .B0(ssrms0_out[15]), 
        .B1(n4811), .Y(n3971) );
  AOI22X1TS U4550 ( .A0(rege_out[1]), .A1(n3980), .B0(n3971), .B1(n4810), .Y(
        n4010) );
  AOI22X1TS U4551 ( .A0(rege_out[2]), .A1(n4111), .B0(n4010), .B1(n4812), .Y(
        n4067) );
  AOI22X1TS U4552 ( .A0(rege_out[3]), .A1(n4235), .B0(n4067), .B1(n4772), .Y(
        n4172) );
  AOI22X1TS U4553 ( .A0(n4293), .A1(aluone_out[31]), .B0(n4044), .B1(n4172), 
        .Y(n3750) );
  OAI31X1TS U4554 ( .A0(n4772), .A1(n4209), .A2(n4070), .B0(n3750), .Y(n3754)
         );
  INVX2TS U4555 ( .A(ssrms0_out[30]), .Y(n3968) );
  NAND3XLTS U4556 ( .A(ssr_ms0[1]), .B(n4418), .C(n3751), .Y(n4117) );
  INVX2TS U4557 ( .A(n4126), .Y(n4298) );
  AOI22X1TS U4558 ( .A0(n4290), .A1(mult1_out[31]), .B0(n4298), .B1(
        ssrms0_out[32]), .Y(n3752) );
  OAI211XLTS U4559 ( .A0(n3968), .A1(n4117), .B0(n3752), .C0(n4135), .Y(n3753)
         );
  OAI21XLTS U4560 ( .A0(n3754), .A1(n3753), .B0(n3756), .Y(n3755) );
  OAI21XLTS U4561 ( .A0(n3756), .A1(n3959), .B0(n3755), .Y(n1910) );
  INVX2TS U4562 ( .A(srmp_out[61]), .Y(n3770) );
  NAND2X1TS U4563 ( .A(sr_mp[1]), .B(n3757), .Y(n3768) );
  AOI22X1TS U4564 ( .A0(n1985), .A1(srmp_out[60]), .B0(n4407), .B1(
        srmp_out[59]), .Y(n3758) );
  NAND2X1TS U4565 ( .A(mult2_out[63]), .B(n4413), .Y(n4305) );
  OAI211XLTS U4566 ( .A0(n3770), .A1(n3764), .B0(n3758), .C0(n4305), .Y(n1875)
         );
  INVX2TS U4567 ( .A(srmp_out[57]), .Y(n3762) );
  AOI22X1TS U4568 ( .A0(n1985), .A1(srmp_out[56]), .B0(n4407), .B1(
        srmp_out[55]), .Y(n3759) );
  OAI211XLTS U4569 ( .A0(n3764), .A1(n3762), .B0(n3759), .C0(n4305), .Y(n1871)
         );
  INVX2TS U4570 ( .A(srmp_out[59]), .Y(n3766) );
  AOI22X1TS U4571 ( .A0(n1985), .A1(srmp_out[58]), .B0(n4407), .B1(
        srmp_out[57]), .Y(n3760) );
  OAI211XLTS U4572 ( .A0(n3764), .A1(n3766), .B0(n3760), .C0(n4305), .Y(n1873)
         );
  AOI22X1TS U4573 ( .A0(n4407), .A1(srmp_out[56]), .B0(n4412), .B1(
        srmp_out[58]), .Y(n3761) );
  OAI211XLTS U4574 ( .A0(n4304), .A1(n3762), .B0(n3761), .C0(n4305), .Y(n1872)
         );
  INVX2TS U4575 ( .A(srmp_out[55]), .Y(n3772) );
  AOI22X1TS U4576 ( .A0(n1985), .A1(srmp_out[54]), .B0(n4407), .B1(
        srmp_out[53]), .Y(n3763) );
  OAI211XLTS U4577 ( .A0(n3764), .A1(n3772), .B0(n3763), .C0(n4305), .Y(n1869)
         );
  AOI22X1TS U4578 ( .A0(n4407), .A1(srmp_out[58]), .B0(n4412), .B1(
        srmp_out[60]), .Y(n3765) );
  OAI211XLTS U4579 ( .A0(n4304), .A1(n3766), .B0(n3765), .C0(n4305), .Y(n1874)
         );
  AOI22X1TS U4580 ( .A0(n1985), .A1(srmp_out[62]), .B0(n4412), .B1(
        srmp_out[63]), .Y(n3767) );
  OAI211XLTS U4581 ( .A0(n3768), .A1(n3770), .B0(n3767), .C0(n4305), .Y(n1877)
         );
  AOI22X1TS U4582 ( .A0(n4407), .A1(srmp_out[60]), .B0(srmp_out[62]), .B1(
        n4412), .Y(n3769) );
  OAI211XLTS U4583 ( .A0(n4304), .A1(n3770), .B0(n3769), .C0(n4305), .Y(n1876)
         );
  AOI22X1TS U4584 ( .A0(n4407), .A1(srmp_out[54]), .B0(n4412), .B1(
        srmp_out[56]), .Y(n3771) );
  OAI211XLTS U4585 ( .A0(n4304), .A1(n3772), .B0(n3771), .C0(n4305), .Y(n1870)
         );
  OR2X1TS U4586 ( .A(sr_mq[1]), .B(sr_mq[0]), .Y(n4484) );
  INVX2TS U4587 ( .A(srmq_out[55]), .Y(n3787) );
  INVX2TS U4588 ( .A(sr_mq[0]), .Y(n3773) );
  NAND2X1TS U4589 ( .A(sr_mq[1]), .B(n3773), .Y(n3780) );
  NAND2X1TS U4590 ( .A(sr_mq[1]), .B(sr_mq[0]), .Y(n3788) );
  AOI22X1TS U4591 ( .A0(n4592), .A1(srmq_out[54]), .B0(n4597), .B1(
        srmq_out[56]), .Y(n3774) );
  NOR2X1TS U4592 ( .A(sr_mq[1]), .B(n3773), .Y(n4515) );
  NAND2X1TS U4593 ( .A(mult2_out[63]), .B(n4595), .Y(n4485) );
  OAI211XLTS U4594 ( .A0(n4484), .A1(n3787), .B0(n3774), .C0(n4485), .Y(n1774)
         );
  INVX2TS U4595 ( .A(srmq_out[61]), .Y(n3782) );
  AOI22X1TS U4596 ( .A0(n1987), .A1(srmq_out[60]), .B0(n4592), .B1(
        srmq_out[59]), .Y(n3775) );
  OAI211XLTS U4597 ( .A0(n3782), .A1(n3788), .B0(n3775), .C0(n4485), .Y(n1779)
         );
  INVX2TS U4598 ( .A(srmq_out[59]), .Y(n3778) );
  AOI22X1TS U4599 ( .A0(n1987), .A1(srmq_out[58]), .B0(n4592), .B1(
        srmq_out[57]), .Y(n3776) );
  OAI211XLTS U4600 ( .A0(n3788), .A1(n3778), .B0(n3776), .C0(n4485), .Y(n1777)
         );
  AOI22X1TS U4601 ( .A0(n4592), .A1(srmq_out[58]), .B0(n4597), .B1(
        srmq_out[60]), .Y(n3777) );
  OAI211XLTS U4602 ( .A0(n4484), .A1(n3778), .B0(n3777), .C0(n4485), .Y(n1778)
         );
  AOI22X1TS U4603 ( .A0(n1987), .A1(srmq_out[62]), .B0(n4597), .B1(
        srmq_out[63]), .Y(n3779) );
  OAI211XLTS U4604 ( .A0(n3780), .A1(n3782), .B0(n3779), .C0(n4485), .Y(n1781)
         );
  AOI22X1TS U4605 ( .A0(n4592), .A1(srmq_out[60]), .B0(srmq_out[62]), .B1(
        n4597), .Y(n3781) );
  OAI211XLTS U4606 ( .A0(n4484), .A1(n3782), .B0(n3781), .C0(n4485), .Y(n1780)
         );
  INVX2TS U4607 ( .A(srmq_out[57]), .Y(n3785) );
  AOI22X1TS U4608 ( .A0(n4592), .A1(srmq_out[56]), .B0(n4597), .B1(
        srmq_out[58]), .Y(n3783) );
  OAI211XLTS U4609 ( .A0(n4484), .A1(n3785), .B0(n3783), .C0(n4485), .Y(n1776)
         );
  AOI22X1TS U4610 ( .A0(n1987), .A1(srmq_out[56]), .B0(n4592), .B1(
        srmq_out[55]), .Y(n3784) );
  OAI211XLTS U4611 ( .A0(n3788), .A1(n3785), .B0(n3784), .C0(n4485), .Y(n1775)
         );
  AOI22X1TS U4612 ( .A0(n1987), .A1(srmq_out[54]), .B0(n4592), .B1(
        srmq_out[53]), .Y(n3786) );
  OAI211XLTS U4613 ( .A0(n3788), .A1(n3787), .B0(n3786), .C0(n4485), .Y(n1773)
         );
  AOI211XLTS U4614 ( .A0(n3812), .A1(n3810), .B0(ssrms0_out[23]), .C0(n3789), 
        .Y(pe_out[3]) );
  AOI21X1TS U4615 ( .A0(n3812), .A1(n4204), .B0(n3790), .Y(n3792) );
  NOR3XLTS U4616 ( .A(ssrms0_out[20]), .B(ssrms0_out[21]), .C(ssrms0_out[22]), 
        .Y(n3791) );
  OAI31X1TS U4617 ( .A0(n3794), .A1(n3793), .A2(n3792), .B0(n3791), .Y(n3795)
         );
  NOR2XLTS U4618 ( .A(ssrms0_out[23]), .B(n3795), .Y(pe_out[2]) );
  INVX2TS U4619 ( .A(n3798), .Y(n3796) );
  AOI22X1TS U4620 ( .A0(n3796), .A1(n3932), .B0(n4819), .B1(count_out[0]), .Y(
        \count/N29 ) );
  OA22X1TS U4621 ( .A0(\C43/DATA3_1 ), .A1(n3799), .B0(count_out[1]), .B1(
        n3798), .Y(\count/N30 ) );
  OAI2BB2XLTS U4622 ( .B0(n3798), .B1(n4075), .A0N(n4819), .A1N(\C43/DATA3_3 ), 
        .Y(\count/N32 ) );
  XOR2XLTS U4623 ( .A(\DP_OP_117J3_124_765/n2 ), .B(count_out[5]), .Y(n3797)
         );
  INVX2TS U4624 ( .A(count_out[5]), .Y(n3881) );
  OAI22X1TS U4625 ( .A0(n3797), .A1(n3799), .B0(n3881), .B1(n3798), .Y(
        \count/N34 ) );
  OA22X1TS U4626 ( .A0(\C43/DATA3_2 ), .A1(n3799), .B0(count_out[2]), .B1(
        n3798), .Y(n4780) );
  NOR4XLTS U4629 ( .A(regsum_out[4]), .B(regsum_out[5]), .C(regsum_out[6]), 
        .D(regsum_out[7]), .Y(n3809) );
  NOR4XLTS U4630 ( .A(regsum_out[0]), .B(regsum_out[1]), .C(regsum_out[2]), 
        .D(regsum_out[3]), .Y(n3808) );
  NOR4XLTS U4631 ( .A(regsum_out[29]), .B(regsum_out[28]), .C(regsum_out[27]), 
        .D(regsum_out[26]), .Y(n3800) );
  NAND3XLTS U4632 ( .A(n3800), .B(n4781), .C(n4775), .Y(n3806) );
  NOR4XLTS U4633 ( .A(regsum_out[12]), .B(regsum_out[13]), .C(regsum_out[14]), 
        .D(regsum_out[15]), .Y(n3804) );
  NOR4XLTS U4634 ( .A(regsum_out[8]), .B(regsum_out[9]), .C(regsum_out[10]), 
        .D(regsum_out[11]), .Y(n3803) );
  NOR4XLTS U4635 ( .A(regsum_out[23]), .B(regsum_out[20]), .C(regsum_out[21]), 
        .D(regsum_out[22]), .Y(n3802) );
  NOR4XLTS U4636 ( .A(regsum_out[16]), .B(regsum_out[17]), .C(regsum_out[18]), 
        .D(regsum_out[19]), .Y(n3801) );
  NAND4XLTS U4637 ( .A(n3804), .B(n3803), .C(n3802), .D(n3801), .Y(n3805) );
  NOR4XLTS U4638 ( .A(regsum_out[30]), .B(regsum_out[31]), .C(n3806), .D(n3805), .Y(n3807) );
  NAND3XLTS U4639 ( .A(n3809), .B(n3808), .C(n3807), .Y(sumorrr_out) );
  INVX2TS U4640 ( .A(ssrms0_out[23]), .Y(n4079) );
  AND4X1TS U4641 ( .A(n3812), .B(n3811), .C(n3810), .D(n4079), .Y(pe_out[4])
         );
  AOI22X1TS U4642 ( .A0(n4290), .A1(mult1_out[63]), .B0(n4274), .B1(
        ssrms0_out[62]), .Y(n3816) );
  NOR3XLTS U4643 ( .A(n3880), .B(n3881), .C(n3813), .Y(n3846) );
  AOI21X1TS U4644 ( .A0(count_out[3]), .A1(n3846), .B0(n4170), .Y(n3843) );
  NOR2XLTS U4645 ( .A(n4234), .B(n3843), .Y(n3815) );
  INVX2TS U4646 ( .A(ssrms0_out[63]), .Y(n3818) );
  INVX2TS U4647 ( .A(n3815), .Y(n3814) );
  AOI32X1TS U4648 ( .A0(n3816), .A1(n3815), .A2(n4135), .B0(n3818), .B1(n3814), 
        .Y(n1942) );
  AOI22X1TS U4649 ( .A0(n4290), .A1(mult1_out[62]), .B0(n4274), .B1(
        ssrms0_out[61]), .Y(n3817) );
  OAI211XLTS U4650 ( .A0(n4126), .A1(n3818), .B0(n3817), .C0(n4135), .Y(n3820)
         );
  AOI31XLTS U4651 ( .A0(count_out[2]), .A1(count_out[1]), .A2(n3932), .B0(
        n3880), .Y(n4243) );
  NOR2XLTS U4652 ( .A(n4243), .B(n3843), .Y(n3819) );
  MX2X1TS U4653 ( .A(ssrms0_out[62]), .B(n3820), .S0(n3819), .Y(n1941) );
  AOI22X1TS U4654 ( .A0(n4290), .A1(mult1_out[61]), .B0(n4274), .B1(
        ssrms0_out[60]), .Y(n3824) );
  AOI31XLTS U4655 ( .A0(count_out[2]), .A1(count_out[0]), .A2(n3931), .B0(
        n3880), .Y(n4252) );
  NOR2XLTS U4656 ( .A(n4252), .B(n3843), .Y(n3823) );
  INVX2TS U4657 ( .A(n4135), .Y(n4297) );
  AOI21X1TS U4658 ( .A0(n4298), .A1(ssrms0_out[62]), .B0(n4297), .Y(n3822) );
  INVX2TS U4659 ( .A(ssrms0_out[61]), .Y(n3826) );
  INVX2TS U4660 ( .A(n3823), .Y(n3821) );
  AOI32X1TS U4661 ( .A0(n3824), .A1(n3823), .A2(n3822), .B0(n3826), .B1(n3821), 
        .Y(n1940) );
  AOI22X1TS U4662 ( .A0(n4290), .A1(mult1_out[60]), .B0(n4274), .B1(
        ssrms0_out[59]), .Y(n3825) );
  OAI211XLTS U4663 ( .A0(n4126), .A1(n3826), .B0(n3825), .C0(n4135), .Y(n3828)
         );
  AOI31XLTS U4664 ( .A0(count_out[2]), .A1(n3932), .A2(n3931), .B0(n3880), .Y(
        n4261) );
  NOR2XLTS U4665 ( .A(n4261), .B(n3843), .Y(n3827) );
  MX2X1TS U4666 ( .A(ssrms0_out[60]), .B(n3828), .S0(n3827), .Y(n1939) );
  AOI22X1TS U4667 ( .A0(n4290), .A1(mult1_out[59]), .B0(n4298), .B1(
        ssrms0_out[60]), .Y(n3832) );
  NOR3XLTS U4668 ( .A(count_out[2]), .B(n3932), .C(n3931), .Y(n3939) );
  NOR2XLTS U4669 ( .A(n3939), .B(n3880), .Y(n4270) );
  NOR2XLTS U4670 ( .A(n4270), .B(n3843), .Y(n3831) );
  AOI21X1TS U4671 ( .A0(n4274), .A1(ssrms0_out[58]), .B0(n4297), .Y(n3830) );
  INVX2TS U4672 ( .A(ssrms0_out[59]), .Y(n3834) );
  INVX2TS U4673 ( .A(n3831), .Y(n3829) );
  AOI32X1TS U4674 ( .A0(n3832), .A1(n3831), .A2(n3830), .B0(n3834), .B1(n3829), 
        .Y(n1938) );
  AOI22X1TS U4675 ( .A0(n4290), .A1(mult1_out[58]), .B0(n4274), .B1(
        ssrms0_out[57]), .Y(n3833) );
  OAI211XLTS U4676 ( .A0(n4126), .A1(n3834), .B0(n3833), .C0(n4135), .Y(n3836)
         );
  NOR3XLTS U4677 ( .A(count_out[0]), .B(count_out[2]), .C(n3931), .Y(n3943) );
  NOR2XLTS U4678 ( .A(n3943), .B(n3880), .Y(n4280) );
  NOR2XLTS U4679 ( .A(n4280), .B(n3843), .Y(n3835) );
  MX2X1TS U4680 ( .A(ssrms0_out[58]), .B(n3836), .S0(n3835), .Y(n1937) );
  AOI22X1TS U4681 ( .A0(n4274), .A1(ssrms0_out[56]), .B0(n4298), .B1(
        ssrms0_out[58]), .Y(n3840) );
  NOR3XLTS U4682 ( .A(count_out[2]), .B(count_out[1]), .C(n3932), .Y(n3949) );
  NOR2XLTS U4683 ( .A(n3949), .B(n3880), .Y(n4292) );
  NOR2XLTS U4684 ( .A(n4292), .B(n3843), .Y(n3839) );
  AOI21X1TS U4685 ( .A0(n4290), .A1(mult1_out[57]), .B0(n4297), .Y(n3838) );
  INVX2TS U4686 ( .A(ssrms0_out[57]), .Y(n3842) );
  INVX2TS U4687 ( .A(n3839), .Y(n3837) );
  AOI32X1TS U4688 ( .A0(n3840), .A1(n3839), .A2(n3838), .B0(n3842), .B1(n3837), 
        .Y(n1936) );
  AOI22X1TS U4689 ( .A0(n4290), .A1(mult1_out[56]), .B0(n4274), .B1(
        ssrms0_out[55]), .Y(n3841) );
  OAI211XLTS U4690 ( .A0(n4126), .A1(n3842), .B0(n3841), .C0(n4135), .Y(n3845)
         );
  NOR2XLTS U4691 ( .A(n4225), .B(n3843), .Y(n3844) );
  MX2X1TS U4692 ( .A(ssrms0_out[56]), .B(n3845), .S0(n3844), .Y(n1935) );
  AOI22X1TS U4693 ( .A0(n4290), .A1(mult1_out[55]), .B0(n4298), .B1(
        ssrms0_out[56]), .Y(n3850) );
  AOI21X1TS U4694 ( .A0(n3846), .A1(n4075), .B0(n4170), .Y(n3877) );
  NOR2XLTS U4695 ( .A(n4234), .B(n3877), .Y(n3849) );
  AOI21X1TS U4696 ( .A0(n4274), .A1(ssrms0_out[54]), .B0(n4297), .Y(n3848) );
  INVX2TS U4697 ( .A(ssrms0_out[55]), .Y(n3852) );
  INVX2TS U4698 ( .A(n3849), .Y(n3847) );
  AOI32X1TS U4699 ( .A0(n3850), .A1(n3849), .A2(n3848), .B0(n3852), .B1(n3847), 
        .Y(n1934) );
  AOI22X1TS U4700 ( .A0(n4290), .A1(mult1_out[54]), .B0(n4274), .B1(
        ssrms0_out[53]), .Y(n3851) );
  OAI211XLTS U4701 ( .A0(n4126), .A1(n3852), .B0(n3851), .C0(n4135), .Y(n3854)
         );
  NOR2XLTS U4702 ( .A(n4243), .B(n3877), .Y(n3853) );
  MX2X1TS U4703 ( .A(ssrms0_out[54]), .B(n3854), .S0(n3853), .Y(n1933) );
  AOI22X1TS U4704 ( .A0(n4274), .A1(ssrms0_out[52]), .B0(n4298), .B1(
        ssrms0_out[54]), .Y(n3858) );
  NOR2XLTS U4705 ( .A(n4252), .B(n3877), .Y(n3857) );
  AOI21X1TS U4706 ( .A0(n4290), .A1(mult1_out[53]), .B0(n4297), .Y(n3856) );
  INVX2TS U4707 ( .A(ssrms0_out[53]), .Y(n3860) );
  INVX2TS U4708 ( .A(n3857), .Y(n3855) );
  AOI32X1TS U4709 ( .A0(n3858), .A1(n3857), .A2(n3856), .B0(n3860), .B1(n3855), 
        .Y(n1932) );
  AOI22X1TS U4710 ( .A0(n4290), .A1(mult1_out[52]), .B0(n4274), .B1(
        ssrms0_out[51]), .Y(n3859) );
  OAI211XLTS U4711 ( .A0(n4126), .A1(n3860), .B0(n3859), .C0(n4135), .Y(n3862)
         );
  NOR2XLTS U4712 ( .A(n4261), .B(n3877), .Y(n3861) );
  MX2X1TS U4713 ( .A(ssrms0_out[52]), .B(n3862), .S0(n3861), .Y(n1931) );
  AOI22X1TS U4714 ( .A0(n4274), .A1(ssrms0_out[50]), .B0(n4298), .B1(
        ssrms0_out[52]), .Y(n3866) );
  NOR2XLTS U4715 ( .A(n4270), .B(n3877), .Y(n3865) );
  AOI21X1TS U4716 ( .A0(n4290), .A1(mult1_out[51]), .B0(n4297), .Y(n3864) );
  INVX2TS U4717 ( .A(ssrms0_out[51]), .Y(n3868) );
  INVX2TS U4718 ( .A(n3865), .Y(n3863) );
  AOI32X1TS U4719 ( .A0(n3866), .A1(n3865), .A2(n3864), .B0(n3868), .B1(n3863), 
        .Y(n1930) );
  AOI22X1TS U4720 ( .A0(n4290), .A1(mult1_out[50]), .B0(n4274), .B1(
        ssrms0_out[49]), .Y(n3867) );
  OAI211XLTS U4721 ( .A0(n4126), .A1(n3868), .B0(n3867), .C0(n4135), .Y(n3870)
         );
  NOR2XLTS U4722 ( .A(n4280), .B(n3877), .Y(n3869) );
  MX2X1TS U4723 ( .A(ssrms0_out[50]), .B(n3870), .S0(n3869), .Y(n1929) );
  AOI22X1TS U4724 ( .A0(n4290), .A1(mult1_out[49]), .B0(n4274), .B1(
        ssrms0_out[48]), .Y(n3874) );
  NOR2XLTS U4725 ( .A(n4292), .B(n3877), .Y(n3873) );
  AOI21X1TS U4726 ( .A0(n4298), .A1(ssrms0_out[50]), .B0(n4297), .Y(n3872) );
  INVX2TS U4727 ( .A(ssrms0_out[49]), .Y(n3876) );
  INVX2TS U4728 ( .A(n3873), .Y(n3871) );
  AOI32X1TS U4729 ( .A0(n3874), .A1(n3873), .A2(n3872), .B0(n3876), .B1(n3871), 
        .Y(n1928) );
  AOI22X1TS U4730 ( .A0(n4290), .A1(mult1_out[48]), .B0(n4274), .B1(
        ssrms0_out[47]), .Y(n3875) );
  OAI211XLTS U4731 ( .A0(n4126), .A1(n3876), .B0(n3875), .C0(n4135), .Y(n3879)
         );
  NOR2XLTS U4732 ( .A(n4225), .B(n3877), .Y(n3878) );
  MX2X1TS U4733 ( .A(ssrms0_out[48]), .B(n3879), .S0(n3878), .Y(n1927) );
  AOI22X1TS U4734 ( .A0(n4290), .A1(mult1_out[47]), .B0(n4298), .B1(
        ssrms0_out[48]), .Y(n3885) );
  NOR3XLTS U4735 ( .A(count_out[4]), .B(n3881), .C(n3880), .Y(n3918) );
  AOI21X1TS U4736 ( .A0(count_out[3]), .A1(n3918), .B0(n4170), .Y(n3911) );
  NOR2XLTS U4737 ( .A(n4234), .B(n3911), .Y(n3884) );
  AOI21X1TS U4738 ( .A0(n4274), .A1(ssrms0_out[46]), .B0(n4297), .Y(n3883) );
  INVX2TS U4739 ( .A(ssrms0_out[47]), .Y(n3887) );
  INVX2TS U4740 ( .A(n3884), .Y(n3882) );
  AOI32X1TS U4741 ( .A0(n3885), .A1(n3884), .A2(n3883), .B0(n3887), .B1(n3882), 
        .Y(n1926) );
  AOI22X1TS U4742 ( .A0(n4290), .A1(mult1_out[46]), .B0(n4274), .B1(
        ssrms0_out[45]), .Y(n3886) );
  OAI211XLTS U4743 ( .A0(n4126), .A1(n3887), .B0(n3886), .C0(n4135), .Y(n3889)
         );
  NOR2XLTS U4744 ( .A(n4243), .B(n3911), .Y(n3888) );
  MX2X1TS U4745 ( .A(ssrms0_out[46]), .B(n3889), .S0(n3888), .Y(n1925) );
  AOI22X1TS U4746 ( .A0(n4274), .A1(ssrms0_out[44]), .B0(n4298), .B1(
        ssrms0_out[46]), .Y(n3893) );
  NOR2XLTS U4747 ( .A(n4252), .B(n3911), .Y(n3892) );
  AOI21X1TS U4748 ( .A0(n4290), .A1(mult1_out[45]), .B0(n4297), .Y(n3891) );
  INVX2TS U4749 ( .A(ssrms0_out[45]), .Y(n3895) );
  INVX2TS U4750 ( .A(n3892), .Y(n3890) );
  AOI32X1TS U4751 ( .A0(n3893), .A1(n3892), .A2(n3891), .B0(n3895), .B1(n3890), 
        .Y(n1924) );
  AOI22X1TS U4752 ( .A0(n4290), .A1(mult1_out[44]), .B0(n4274), .B1(
        ssrms0_out[43]), .Y(n3894) );
  OAI211XLTS U4753 ( .A0(n4126), .A1(n3895), .B0(n3894), .C0(n4135), .Y(n3897)
         );
  NOR2XLTS U4754 ( .A(n4261), .B(n3911), .Y(n3896) );
  MX2X1TS U4755 ( .A(ssrms0_out[44]), .B(n3897), .S0(n3896), .Y(n1923) );
  AOI22X1TS U4756 ( .A0(n4290), .A1(mult1_out[43]), .B0(n4274), .B1(
        ssrms0_out[42]), .Y(n3901) );
  NOR2XLTS U4757 ( .A(n4270), .B(n3911), .Y(n3900) );
  AOI21X1TS U4758 ( .A0(n4298), .A1(ssrms0_out[44]), .B0(n4297), .Y(n3899) );
  INVX2TS U4759 ( .A(ssrms0_out[43]), .Y(n3903) );
  INVX2TS U4760 ( .A(n3900), .Y(n3898) );
  AOI32X1TS U4761 ( .A0(n3901), .A1(n3900), .A2(n3899), .B0(n3903), .B1(n3898), 
        .Y(n1922) );
  AOI22X1TS U4762 ( .A0(n4290), .A1(mult1_out[42]), .B0(n4274), .B1(
        ssrms0_out[41]), .Y(n3902) );
  OAI211XLTS U4763 ( .A0(n4126), .A1(n3903), .B0(n3902), .C0(n4135), .Y(n3905)
         );
  INVX2TS U4764 ( .A(n3911), .Y(n3907) );
  OAI21XLTS U4765 ( .A0(n4170), .A1(n3943), .B0(n3907), .Y(n3904) );
  MX2X1TS U4766 ( .A(n3905), .B(ssrms0_out[42]), .S0(n3904), .Y(n1921) );
  AO22XLTS U4767 ( .A0(n4274), .A1(ssrms0_out[40]), .B0(n4298), .B1(
        ssrms0_out[42]), .Y(n3906) );
  AOI211XLTS U4768 ( .A0(n4290), .A1(mult1_out[41]), .B0(n4297), .C0(n3906), 
        .Y(n3910) );
  INVX2TS U4769 ( .A(ssrms0_out[41]), .Y(n3909) );
  OAI21XLTS U4770 ( .A0(n4170), .A1(n3949), .B0(n3907), .Y(n3908) );
  MXI2XLTS U4771 ( .A(n3910), .B(n3909), .S0(n3908), .Y(n1920) );
  AOI22X1TS U4772 ( .A0(n4290), .A1(mult1_out[40]), .B0(n4298), .B1(
        ssrms0_out[41]), .Y(n3915) );
  NOR2XLTS U4773 ( .A(n4225), .B(n3911), .Y(n3914) );
  AOI21X1TS U4774 ( .A0(n4274), .A1(ssrms0_out[39]), .B0(n4297), .Y(n3913) );
  INVX2TS U4775 ( .A(ssrms0_out[40]), .Y(n3917) );
  INVX2TS U4776 ( .A(n3914), .Y(n3912) );
  AOI32X1TS U4777 ( .A0(n3915), .A1(n3914), .A2(n3913), .B0(n3917), .B1(n3912), 
        .Y(n1919) );
  AOI22X1TS U4778 ( .A0(n4290), .A1(mult1_out[39]), .B0(n4274), .B1(
        ssrms0_out[38]), .Y(n3916) );
  OAI211XLTS U4779 ( .A0(n4126), .A1(n3917), .B0(n3916), .C0(n4135), .Y(n3920)
         );
  AOI21X1TS U4780 ( .A0(n3918), .A1(n4075), .B0(n4170), .Y(n3952) );
  NOR2XLTS U4781 ( .A(n4234), .B(n3952), .Y(n3919) );
  MX2X1TS U4782 ( .A(ssrms0_out[39]), .B(n3920), .S0(n3919), .Y(n1918) );
  INVX2TS U4783 ( .A(ssrms0_out[38]), .Y(n3926) );
  AO22XLTS U4784 ( .A0(n4274), .A1(ssrms0_out[37]), .B0(n4298), .B1(
        ssrms0_out[39]), .Y(n3921) );
  AOI211XLTS U4785 ( .A0(n4290), .A1(mult1_out[38]), .B0(n4297), .C0(n3921), 
        .Y(n3924) );
  NAND3XLTS U4786 ( .A(count_out[2]), .B(count_out[1]), .C(n3932), .Y(n3922)
         );
  AOI21X1TS U4787 ( .A0(n3934), .A1(n3922), .B0(n3952), .Y(n3923) );
  MXI2XLTS U4788 ( .A(n3926), .B(n3924), .S0(n3923), .Y(n1917) );
  AOI22X1TS U4789 ( .A0(n4290), .A1(mult1_out[37]), .B0(n4274), .B1(
        ssrms0_out[36]), .Y(n3925) );
  OAI211XLTS U4790 ( .A0(n4126), .A1(n3926), .B0(n3925), .C0(n4135), .Y(n3929)
         );
  NAND3XLTS U4791 ( .A(count_out[2]), .B(count_out[0]), .C(n3931), .Y(n3927)
         );
  AOI21X1TS U4792 ( .A0(n3934), .A1(n3927), .B0(n3952), .Y(n3928) );
  MX2X1TS U4793 ( .A(ssrms0_out[37]), .B(n3929), .S0(n3928), .Y(n1916) );
  INVX2TS U4794 ( .A(ssrms0_out[36]), .Y(n3938) );
  AO22XLTS U4795 ( .A0(n4274), .A1(ssrms0_out[35]), .B0(n4298), .B1(
        ssrms0_out[37]), .Y(n3930) );
  AOI211XLTS U4796 ( .A0(n4290), .A1(mult1_out[36]), .B0(n4297), .C0(n3930), 
        .Y(n3936) );
  NAND3XLTS U4797 ( .A(count_out[2]), .B(n3932), .C(n3931), .Y(n3933) );
  AOI21X1TS U4798 ( .A0(n3934), .A1(n3933), .B0(n3952), .Y(n3935) );
  MXI2XLTS U4799 ( .A(n3938), .B(n3936), .S0(n3935), .Y(n1915) );
  AOI22X1TS U4800 ( .A0(n4290), .A1(mult1_out[35]), .B0(n4274), .B1(
        ssrms0_out[34]), .Y(n3937) );
  OAI211XLTS U4801 ( .A0(n4126), .A1(n3938), .B0(n3937), .C0(n4135), .Y(n3941)
         );
  INVX2TS U4802 ( .A(n3952), .Y(n3948) );
  OAI21XLTS U4803 ( .A0(n4170), .A1(n3939), .B0(n3948), .Y(n3940) );
  MX2X1TS U4804 ( .A(n3941), .B(ssrms0_out[35]), .S0(n3940), .Y(n1914) );
  AO22XLTS U4805 ( .A0(n4274), .A1(ssrms0_out[33]), .B0(n4298), .B1(
        ssrms0_out[35]), .Y(n3942) );
  AOI211XLTS U4806 ( .A0(n4290), .A1(mult1_out[34]), .B0(n4297), .C0(n3942), 
        .Y(n3945) );
  INVX2TS U4807 ( .A(ssrms0_out[34]), .Y(n3947) );
  OAI21XLTS U4808 ( .A0(n4170), .A1(n3943), .B0(n3948), .Y(n3944) );
  MXI2XLTS U4809 ( .A(n3945), .B(n3947), .S0(n3944), .Y(n1913) );
  AOI22X1TS U4810 ( .A0(n4290), .A1(mult1_out[33]), .B0(n4274), .B1(
        ssrms0_out[32]), .Y(n3946) );
  OAI211XLTS U4811 ( .A0(n4126), .A1(n3947), .B0(n3946), .C0(n4135), .Y(n3951)
         );
  OAI21XLTS U4812 ( .A0(n4170), .A1(n3949), .B0(n3948), .Y(n3950) );
  MX2X1TS U4813 ( .A(n3951), .B(ssrms0_out[33]), .S0(n3950), .Y(n1912) );
  AOI22X1TS U4814 ( .A0(n4290), .A1(mult1_out[32]), .B0(n4298), .B1(
        ssrms0_out[33]), .Y(n3957) );
  NOR2XLTS U4815 ( .A(n4225), .B(n3952), .Y(n3956) );
  AOI21X1TS U4816 ( .A0(ssrms0_out[31]), .A1(n4274), .B0(n4297), .Y(n3955) );
  INVX2TS U4817 ( .A(ssrms0_out[32]), .Y(n3954) );
  INVX2TS U4818 ( .A(n3956), .Y(n3953) );
  AOI32X1TS U4819 ( .A0(n3957), .A1(n3956), .A2(n3955), .B0(n3954), .B1(n3953), 
        .Y(n1911) );
  AOI22X1TS U4820 ( .A0(ssrms0_out[29]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[30]), .Y(n3958) );
  OAI211XLTS U4821 ( .A0(n3959), .A1(n4126), .B0(n3958), .C0(n4135), .Y(n3960)
         );
  AOI21X1TS U4822 ( .A0(n4293), .A1(aluone_out[30]), .B0(n3960), .Y(n3966) );
  NOR2XLTS U4823 ( .A(n4050), .B(n4243), .Y(n3965) );
  NAND2X1TS U4824 ( .A(rege_out[3]), .B(n4778), .Y(n4142) );
  AOI22X1TS U4825 ( .A0(rege_out[0]), .A1(ssrms0_out[15]), .B0(ssrms0_out[16]), 
        .B1(n4811), .Y(n3996) );
  AOI22X1TS U4826 ( .A0(rege_out[0]), .A1(ssrms0_out[17]), .B0(ssrms0_out[18]), 
        .B1(n4811), .Y(n3999) );
  AOI22X1TS U4827 ( .A0(rege_out[1]), .A1(n3996), .B0(n3999), .B1(n4810), .Y(
        n4021) );
  AOI22X1TS U4828 ( .A0(rege_out[0]), .A1(ssrms0_out[19]), .B0(ssrms0_out[20]), 
        .B1(n4811), .Y(n3998) );
  AOI22X1TS U4829 ( .A0(rege_out[0]), .A1(ssrms0_out[21]), .B0(ssrms0_out[22]), 
        .B1(n4811), .Y(n4000) );
  AOI22X1TS U4830 ( .A0(rege_out[1]), .A1(n3998), .B0(n4000), .B1(n4810), .Y(
        n4026) );
  AOI22X1TS U4831 ( .A0(rege_out[2]), .A1(n4021), .B0(n4026), .B1(n4812), .Y(
        n4081) );
  NAND2X1TS U4832 ( .A(rege_out[0]), .B(ssrms0_out[23]), .Y(n4023) );
  NOR3XLTS U4833 ( .A(rege_out[3]), .B(rege_out[4]), .C(n4812), .Y(n4058) );
  NAND2X1TS U4834 ( .A(rege_out[1]), .B(n4058), .Y(n3974) );
  OAI22X1TS U4835 ( .A0(n4142), .A1(n4081), .B0(n4023), .B1(n3974), .Y(n3962)
         );
  AOI22X1TS U4836 ( .A0(rege_out[0]), .A1(ssrms0_out[1]), .B0(ssrms0_out[2]), 
        .B1(n4811), .Y(n3988) );
  OAI32X1TS U4837 ( .A0(n4810), .A1(rege_out[0]), .A2(n3961), .B0(rege_out[1]), 
        .B1(n3988), .Y(n4019) );
  AOI22X1TS U4838 ( .A0(rege_out[0]), .A1(ssrms0_out[3]), .B0(ssrms0_out[4]), 
        .B1(n4811), .Y(n3987) );
  AOI22X1TS U4839 ( .A0(rege_out[0]), .A1(ssrms0_out[5]), .B0(ssrms0_out[6]), 
        .B1(n4811), .Y(n3991) );
  AOI22X1TS U4840 ( .A0(rege_out[1]), .A1(n3987), .B0(n3991), .B1(n4810), .Y(
        n4123) );
  AOI22X1TS U4841 ( .A0(rege_out[2]), .A1(n4019), .B0(n4123), .B1(n4812), .Y(
        n4245) );
  AOI22X1TS U4842 ( .A0(rege_out[0]), .A1(ssrms0_out[7]), .B0(ssrms0_out[8]), 
        .B1(n4811), .Y(n3990) );
  AOI22X1TS U4843 ( .A0(rege_out[0]), .A1(ssrms0_out[9]), .B0(ssrms0_out[10]), 
        .B1(n4811), .Y(n3993) );
  AOI22X1TS U4844 ( .A0(rege_out[1]), .A1(n3990), .B0(n3993), .B1(n4810), .Y(
        n4122) );
  AOI22X1TS U4845 ( .A0(rege_out[0]), .A1(ssrms0_out[11]), .B0(ssrms0_out[12]), 
        .B1(n4811), .Y(n3992) );
  AOI22X1TS U4846 ( .A0(rege_out[0]), .A1(ssrms0_out[13]), .B0(ssrms0_out[14]), 
        .B1(n4811), .Y(n3997) );
  AOI22X1TS U4847 ( .A0(rege_out[1]), .A1(n3992), .B0(n3997), .B1(n4810), .Y(
        n4022) );
  AOI22X1TS U4848 ( .A0(rege_out[2]), .A1(n4122), .B0(n4022), .B1(n4812), .Y(
        n4080) );
  AOI22X1TS U4849 ( .A0(rege_out[3]), .A1(n4245), .B0(n4080), .B1(n4772), .Y(
        n4179) );
  AOI22X1TS U4850 ( .A0(n4145), .A1(n3962), .B0(n4044), .B1(n4179), .Y(n3964)
         );
  INVX2TS U4851 ( .A(n3965), .Y(n3963) );
  AOI32X1TS U4852 ( .A0(n3966), .A1(n3965), .A2(n3964), .B0(n3968), .B1(n3963), 
        .Y(n1909) );
  AOI22X1TS U4853 ( .A0(ssrms0_out[28]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[29]), .Y(n3967) );
  OAI211XLTS U4854 ( .A0(n3968), .A1(n4126), .B0(n3967), .C0(n4135), .Y(n3969)
         );
  AOI21X1TS U4855 ( .A0(n4293), .A1(aluone_out[29]), .B0(n3969), .Y(n3986) );
  NOR2XLTS U4856 ( .A(n4050), .B(n4252), .Y(n3985) );
  AOI22X1TS U4857 ( .A0(rege_out[1]), .A1(n3971), .B0(n3970), .B1(n4810), .Y(
        n4035) );
  AOI22X1TS U4858 ( .A0(rege_out[1]), .A1(n3973), .B0(n3972), .B1(n4810), .Y(
        n4037) );
  AOI22X1TS U4859 ( .A0(rege_out[2]), .A1(n4035), .B0(n4037), .B1(n4812), .Y(
        n4092) );
  OAI22X1TS U4860 ( .A0(n4040), .A1(n3974), .B0(n4092), .B1(n4142), .Y(n3982)
         );
  NOR2XLTS U4861 ( .A(rege_out[1]), .B(n3975), .Y(n4042) );
  AOI22X1TS U4862 ( .A0(rege_out[1]), .A1(n3977), .B0(n3976), .B1(n4810), .Y(
        n4140) );
  AOI22X1TS U4863 ( .A0(rege_out[2]), .A1(n4042), .B0(n4140), .B1(n4812), .Y(
        n4254) );
  AOI22X1TS U4864 ( .A0(rege_out[1]), .A1(n3979), .B0(n3978), .B1(n4810), .Y(
        n4139) );
  AOI22X1TS U4865 ( .A0(rege_out[1]), .A1(n3981), .B0(n3980), .B1(n4810), .Y(
        n4036) );
  AOI22X1TS U4866 ( .A0(rege_out[2]), .A1(n4139), .B0(n4036), .B1(n4812), .Y(
        n4089) );
  AOI22X1TS U4867 ( .A0(rege_out[3]), .A1(n4254), .B0(n4089), .B1(n4772), .Y(
        n4186) );
  AOI22X1TS U4868 ( .A0(n4145), .A1(n3982), .B0(n4044), .B1(n4186), .Y(n3984)
         );
  INVX2TS U4869 ( .A(ssrms0_out[29]), .Y(n3995) );
  INVX2TS U4870 ( .A(n3985), .Y(n3983) );
  AOI32X1TS U4871 ( .A0(n3986), .A1(n3985), .A2(n3984), .B0(n3995), .B1(n3983), 
        .Y(n1908) );
  INVX2TS U4872 ( .A(ssrms0_out[28]), .Y(n4008) );
  AOI22X1TS U4873 ( .A0(rege_out[1]), .A1(n3988), .B0(n3987), .B1(n4810), .Y(
        n4153) );
  AOI22X1TS U4874 ( .A0(rege_out[2]), .A1(n3989), .B0(n4153), .B1(n4812), .Y(
        n4263) );
  AOI22X1TS U4875 ( .A0(rege_out[1]), .A1(n3991), .B0(n3990), .B1(n4810), .Y(
        n4154) );
  AOI22X1TS U4876 ( .A0(rege_out[1]), .A1(n3993), .B0(n3992), .B1(n4810), .Y(
        n4055) );
  AOI22X1TS U4877 ( .A0(rege_out[2]), .A1(n4154), .B0(n4055), .B1(n4812), .Y(
        n4102) );
  AOI22X1TS U4878 ( .A0(rege_out[3]), .A1(n4263), .B0(n4102), .B1(n4772), .Y(
        n4193) );
  AOI22X1TS U4879 ( .A0(ssrms0_out[27]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[28]), .Y(n3994) );
  OAI211XLTS U4880 ( .A0(n3995), .A1(n4126), .B0(n3994), .C0(n4135), .Y(n4004)
         );
  INVX2TS U4881 ( .A(n4142), .Y(n4152) );
  AO22XLTS U4882 ( .A0(rege_out[1]), .A1(n3997), .B0(n4810), .B1(n3996), .Y(
        n4056) );
  AOI22X1TS U4883 ( .A0(rege_out[1]), .A1(n3999), .B0(n4810), .B1(n3998), .Y(
        n4057) );
  AOI2BB2XLTS U4884 ( .B0(rege_out[2]), .B1(n4056), .A0N(n4057), .A1N(
        rege_out[2]), .Y(n4103) );
  AOI22X1TS U4885 ( .A0(rege_out[1]), .A1(n4000), .B0(n4023), .B1(n4810), .Y(
        n4051) );
  AOI22X1TS U4886 ( .A0(n4152), .A1(n4103), .B0(n4058), .B1(n4051), .Y(n4002)
         );
  INVX2TS U4887 ( .A(n4293), .Y(n4282) );
  OAI22X1TS U4888 ( .A0(n4002), .A1(n4162), .B0(n4001), .B1(n4282), .Y(n4003)
         );
  AOI211XLTS U4889 ( .A0(n4044), .A1(n4193), .B0(n4004), .C0(n4003), .Y(n4006)
         );
  NOR2XLTS U4890 ( .A(n4050), .B(n4261), .Y(n4005) );
  MXI2XLTS U4891 ( .A(n4008), .B(n4006), .S0(n4005), .Y(n1907) );
  INVX2TS U4892 ( .A(ssrms0_out[27]), .Y(n4029) );
  AOI22X1TS U4893 ( .A0(ssrms0_out[26]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[27]), .Y(n4007) );
  OAI211XLTS U4894 ( .A0(n4008), .A1(n4126), .B0(n4007), .C0(n4135), .Y(n4016)
         );
  AO22XLTS U4895 ( .A0(rege_out[2]), .A1(n4010), .B0(n4812), .B1(n4009), .Y(
        n4112) );
  AOI22X1TS U4896 ( .A0(n4011), .A1(n4058), .B0(n4152), .B1(n4112), .Y(n4014)
         );
  INVX2TS U4897 ( .A(n4044), .Y(n4013) );
  NAND2X1TS U4898 ( .A(n4772), .B(n4812), .Y(n4053) );
  CLKAND2X2TS U4899 ( .A(n4012), .B(n4812), .Y(n4272) );
  OAI222X1TS U4900 ( .A0(n4812), .A1(n4110), .B0(n4053), .B1(n4111), .C0(n4772), .C1(n4272), .Y(n4200) );
  OAI22X1TS U4901 ( .A0(n4014), .A1(n4162), .B0(n4013), .B1(n4200), .Y(n4015)
         );
  AOI211XLTS U4902 ( .A0(n4293), .A1(aluone_out[27]), .B0(n4016), .C0(n4015), 
        .Y(n4018) );
  NOR2XLTS U4903 ( .A(n4050), .B(n4270), .Y(n4017) );
  MXI2XLTS U4904 ( .A(n4029), .B(n4018), .S0(n4017), .Y(n1906) );
  INVX2TS U4905 ( .A(ssrms0_out[26]), .Y(n4034) );
  NAND2X1TS U4906 ( .A(n4812), .B(n4019), .Y(n4281) );
  OAI32X1TS U4907 ( .A0(rege_out[2]), .A1(rege_out[3]), .A2(n4122), .B0(n4123), 
        .B1(n4812), .Y(n4020) );
  AO21XLTS U4908 ( .A0(rege_out[3]), .A1(n4281), .B0(n4020), .Y(n4208) );
  AOI22X1TS U4909 ( .A0(rege_out[2]), .A1(n4022), .B0(n4021), .B1(n4812), .Y(
        n4128) );
  NOR3XLTS U4910 ( .A(rege_out[2]), .B(n4810), .C(n4023), .Y(n4024) );
  AOI2BB2XLTS U4911 ( .B0(n4152), .B1(n4128), .A0N(n4024), .A1N(n4082), .Y(
        n4025) );
  AOI31XLTS U4912 ( .A0(rege_out[2]), .A1(n4026), .A2(n4772), .B0(n4025), .Y(
        n4027) );
  AOI211XLTS U4913 ( .A0(rege_out[4]), .A1(n4208), .B0(n4027), .C0(n4162), .Y(
        n4031) );
  AOI22X1TS U4914 ( .A0(ssrms0_out[25]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[26]), .Y(n4028) );
  OAI211XLTS U4915 ( .A0(n4029), .A1(n4126), .B0(n4028), .C0(n4135), .Y(n4030)
         );
  AOI211XLTS U4916 ( .A0(n4293), .A1(aluone_out[26]), .B0(n4031), .C0(n4030), 
        .Y(n4033) );
  NOR2XLTS U4917 ( .A(n4050), .B(n4280), .Y(n4032) );
  MXI2XLTS U4918 ( .A(n4034), .B(n4033), .S0(n4032), .Y(n1905) );
  AO22XLTS U4919 ( .A0(rege_out[2]), .A1(n4036), .B0(n4812), .B1(n4035), .Y(
        n4143) );
  AOI22X1TS U4920 ( .A0(n4152), .A1(n4143), .B0(n4058), .B1(n4037), .Y(n4047)
         );
  NAND2X1TS U4921 ( .A(rege_out[1]), .B(n4812), .Y(n4039) );
  AOI22X1TS U4922 ( .A0(ssrms0_out[26]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[25]), .Y(n4038) );
  OAI31X1TS U4923 ( .A0(n4040), .A1(n4039), .A2(n4294), .B0(n4038), .Y(n4041)
         );
  AOI211XLTS U4924 ( .A0(ssrms0_out[24]), .A1(n4274), .B0(n4297), .C0(n4041), 
        .Y(n4046) );
  NAND2X1TS U4925 ( .A(n4042), .B(n4812), .Y(n4295) );
  OAI21XLTS U4926 ( .A0(n4140), .A1(n4812), .B0(n4772), .Y(n4043) );
  AOI2BB2XLTS U4927 ( .B0(n4295), .B1(n4043), .A0N(n4139), .A1N(n4053), .Y(
        n4217) );
  AOI22X1TS U4928 ( .A0(n4044), .A1(n4217), .B0(n4293), .B1(aluone_out[25]), 
        .Y(n4045) );
  OAI211XLTS U4929 ( .A0(n4047), .A1(n4162), .B0(n4046), .C0(n4045), .Y(n4049)
         );
  NOR2XLTS U4930 ( .A(n4050), .B(n4292), .Y(n4048) );
  MX2X1TS U4931 ( .A(ssrms0_out[25]), .B(n4049), .S0(n4048), .Y(n1904) );
  AOI22X1TS U4932 ( .A0(ssrms0_out[25]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[24]), .Y(n4066) );
  NOR2XLTS U4933 ( .A(n4050), .B(n4225), .Y(n4065) );
  INVX2TS U4934 ( .A(n4051), .Y(n4052) );
  OAI31X1TS U4935 ( .A0(n4052), .A1(n4209), .A2(n4053), .B0(n4135), .Y(n4062)
         );
  OAI22X1TS U4936 ( .A0(n4153), .A1(n4812), .B0(n4154), .B1(n4053), .Y(n4054)
         );
  AOI21X1TS U4937 ( .A0(rege_out[3]), .A1(n4157), .B0(n4054), .Y(n4226) );
  AOI2BB2XLTS U4938 ( .B0(n4056), .B1(n4812), .A0N(n4812), .A1N(n4055), .Y(
        n4159) );
  AOI222XLTS U4939 ( .A0(rege_out[4]), .A1(n4226), .B0(n4152), .B1(n4159), 
        .C0(n4058), .C1(n4057), .Y(n4060) );
  OAI22X1TS U4940 ( .A0(n4060), .A1(n4162), .B0(n4059), .B1(n4282), .Y(n4061)
         );
  AOI211XLTS U4941 ( .A0(ssrms0_out[23]), .A1(n4274), .B0(n4062), .C0(n4061), 
        .Y(n4064) );
  INVX2TS U4942 ( .A(ssrms0_out[24]), .Y(n4069) );
  INVX2TS U4943 ( .A(n4065), .Y(n4063) );
  AOI32X1TS U4944 ( .A0(n4066), .A1(n4065), .A2(n4064), .B0(n4069), .B1(n4063), 
        .Y(n1903) );
  NAND2X1TS U4945 ( .A(rege_out[4]), .B(n4772), .Y(n4156) );
  OAI22X1TS U4946 ( .A0(n4235), .A1(n4156), .B0(n4067), .B1(n4142), .Y(n4074)
         );
  AOI22X1TS U4947 ( .A0(ssrms0_out[22]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[23]), .Y(n4068) );
  OAI211XLTS U4948 ( .A0(n4069), .A1(n4126), .B0(n4068), .C0(n4135), .Y(n4073)
         );
  OAI22X1TS U4949 ( .A0(n4071), .A1(n4282), .B0(n4070), .B1(n4294), .Y(n4072)
         );
  AOI211XLTS U4950 ( .A0(n4145), .A1(n4074), .B0(n4073), .C0(n4072), .Y(n4078)
         );
  AOI21X1TS U4951 ( .A0(n4076), .A1(n4075), .B0(n4170), .Y(n4151) );
  NOR2XLTS U4952 ( .A(n4234), .B(n4151), .Y(n4077) );
  MXI2XLTS U4953 ( .A(n4079), .B(n4078), .S0(n4077), .Y(n1902) );
  AOI22X1TS U4954 ( .A0(ssrms0_out[21]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[22]), .Y(n4088) );
  NOR2XLTS U4955 ( .A(n4243), .B(n4151), .Y(n4087) );
  OAI222X1TS U4956 ( .A0(n4082), .A1(n4081), .B0(n4156), .B1(n4245), .C0(n4142), .C1(n4080), .Y(n4083) );
  AO22XLTS U4957 ( .A0(n4293), .A1(aluone_out[22]), .B0(n4145), .B1(n4083), 
        .Y(n4084) );
  AOI211XLTS U4958 ( .A0(ssrms0_out[23]), .A1(n4298), .B0(n4297), .C0(n4084), 
        .Y(n4086) );
  INVX2TS U4959 ( .A(n4087), .Y(n4085) );
  AOI32X1TS U4960 ( .A0(n4088), .A1(n4087), .A2(n4086), .B0(n4091), .B1(n4085), 
        .Y(n1901) );
  OAI22X1TS U4961 ( .A0(n4254), .A1(n4156), .B0(n4142), .B1(n4089), .Y(n4096)
         );
  AOI22X1TS U4962 ( .A0(ssrms0_out[20]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[21]), .Y(n4090) );
  OAI211XLTS U4963 ( .A0(n4091), .A1(n4126), .B0(n4090), .C0(n4135), .Y(n4095)
         );
  OAI22X1TS U4964 ( .A0(n4093), .A1(n4282), .B0(n4092), .B1(n4294), .Y(n4094)
         );
  AOI211XLTS U4965 ( .A0(n4145), .A1(n4096), .B0(n4095), .C0(n4094), .Y(n4098)
         );
  NOR2XLTS U4966 ( .A(n4252), .B(n4151), .Y(n4097) );
  MXI2XLTS U4967 ( .A(n4100), .B(n4098), .S0(n4097), .Y(n1900) );
  AOI22X1TS U4968 ( .A0(ssrms0_out[19]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[20]), .Y(n4099) );
  OAI211XLTS U4969 ( .A0(n4100), .A1(n4126), .B0(n4099), .C0(n4135), .Y(n4101)
         );
  AOI21X1TS U4970 ( .A0(n4293), .A1(aluone_out[20]), .B0(n4101), .Y(n4109) );
  NOR2XLTS U4971 ( .A(n4261), .B(n4151), .Y(n4108) );
  OAI22X1TS U4972 ( .A0(n4263), .A1(n4156), .B0(n4142), .B1(n4102), .Y(n4104)
         );
  INVX2TS U4973 ( .A(n4294), .Y(n4271) );
  AOI22X1TS U4974 ( .A0(n4145), .A1(n4104), .B0(n4103), .B1(n4271), .Y(n4107)
         );
  INVX2TS U4975 ( .A(n4108), .Y(n4105) );
  AOI32X1TS U4976 ( .A0(n4109), .A1(n4108), .A2(n4107), .B0(n4106), .B1(n4105), 
        .Y(n1899) );
  OAI221XLTS U4977 ( .A0(rege_out[2]), .A1(n4111), .B0(n4812), .B1(n4110), 
        .C0(n4152), .Y(n4115) );
  INVX2TS U4978 ( .A(n4156), .Y(n4113) );
  AOI22X1TS U4979 ( .A0(n4272), .A1(n4113), .B0(n4112), .B1(n4160), .Y(n4114)
         );
  AOI21X1TS U4980 ( .A0(n4115), .A1(n4114), .B0(n4162), .Y(n4119) );
  AOI22X1TS U4981 ( .A0(ssrms0_out[20]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[19]), .Y(n4116) );
  OAI211XLTS U4982 ( .A0(n4137), .A1(n4117), .B0(n4116), .C0(n4135), .Y(n4118)
         );
  AOI211XLTS U4983 ( .A0(n4293), .A1(aluone_out[19]), .B0(n4119), .C0(n4118), 
        .Y(n4121) );
  NOR2XLTS U4984 ( .A(n4270), .B(n4151), .Y(n4120) );
  MXI2XLTS U4985 ( .A(n4127), .B(n4121), .S0(n4120), .Y(n1898) );
  AOI22X1TS U4986 ( .A0(rege_out[2]), .A1(n4123), .B0(n4122), .B1(n4812), .Y(
        n4124) );
  OAI22X1TS U4987 ( .A0(n4142), .A1(n4124), .B0(n4281), .B1(n4156), .Y(n4132)
         );
  AOI22X1TS U4988 ( .A0(ssrms0_out[17]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[18]), .Y(n4125) );
  OAI211XLTS U4989 ( .A0(n4127), .A1(n4126), .B0(n4125), .C0(n4135), .Y(n4131)
         );
  OAI22X1TS U4990 ( .A0(n4129), .A1(n4282), .B0(n4128), .B1(n4294), .Y(n4130)
         );
  AOI211XLTS U4991 ( .A0(n4145), .A1(n4132), .B0(n4131), .C0(n4130), .Y(n4134)
         );
  NOR2XLTS U4992 ( .A(n4280), .B(n4151), .Y(n4133) );
  MXI2XLTS U4993 ( .A(n4137), .B(n4134), .S0(n4133), .Y(n1897) );
  AOI22X1TS U4994 ( .A0(ssrms0_out[16]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[17]), .Y(n4136) );
  OAI211XLTS U4995 ( .A0(n4137), .A1(n4126), .B0(n4136), .C0(n4135), .Y(n4138)
         );
  AOI21X1TS U4996 ( .A0(n4293), .A1(aluone_out[17]), .B0(n4138), .Y(n4150) );
  NOR2XLTS U4997 ( .A(n4292), .B(n4151), .Y(n4149) );
  AOI22X1TS U4998 ( .A0(rege_out[2]), .A1(n4140), .B0(n4139), .B1(n4812), .Y(
        n4141) );
  OAI22X1TS U4999 ( .A0(n4142), .A1(n4141), .B0(n4295), .B1(n4156), .Y(n4144)
         );
  AOI22X1TS U5000 ( .A0(n4145), .A1(n4144), .B0(n4143), .B1(n4271), .Y(n4148)
         );
  INVX2TS U5001 ( .A(n4149), .Y(n4146) );
  AOI32X1TS U5002 ( .A0(n4150), .A1(n4149), .A2(n4148), .B0(n4147), .B1(n4146), 
        .Y(n1896) );
  AOI22X1TS U5003 ( .A0(ssrms0_out[17]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[16]), .Y(n4169) );
  NOR2XLTS U5004 ( .A(n4225), .B(n4151), .Y(n4168) );
  OAI221XLTS U5005 ( .A0(rege_out[2]), .A1(n4154), .B0(n4812), .B1(n4153), 
        .C0(n4152), .Y(n4155) );
  OAI21XLTS U5006 ( .A0(n4157), .A1(n4156), .B0(n4155), .Y(n4158) );
  AOI21X1TS U5007 ( .A0(n4160), .A1(n4159), .B0(n4158), .Y(n4163) );
  OAI22X1TS U5008 ( .A0(n4163), .A1(n4162), .B0(n4161), .B1(n4282), .Y(n4164)
         );
  AOI211XLTS U5009 ( .A0(ssrms0_out[15]), .A1(n4274), .B0(n4297), .C0(n4164), 
        .Y(n4167) );
  INVX2TS U5010 ( .A(n4168), .Y(n4165) );
  AOI32X1TS U5011 ( .A0(n4169), .A1(n4168), .A2(n4167), .B0(n4166), .B1(n4165), 
        .Y(n1895) );
  AOI22X1TS U5012 ( .A0(ssrms0_out[16]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[15]), .Y(n4178) );
  AOI21X1TS U5013 ( .A0(count_out[3]), .A1(n4171), .B0(n4170), .Y(n4224) );
  NOR2XLTS U5014 ( .A(n4234), .B(n4224), .Y(n4177) );
  INVX2TS U5015 ( .A(n4209), .Y(n4227) );
  AO22XLTS U5016 ( .A0(n4293), .A1(aluone_out[15]), .B0(n4227), .B1(n4172), 
        .Y(n4173) );
  AOI211XLTS U5017 ( .A0(ssrms0_out[14]), .A1(n4274), .B0(n4297), .C0(n4173), 
        .Y(n4176) );
  INVX2TS U5018 ( .A(n4177), .Y(n4174) );
  AOI32X1TS U5019 ( .A0(n4178), .A1(n4177), .A2(n4176), .B0(n4175), .B1(n4174), 
        .Y(n1894) );
  AOI22X1TS U5020 ( .A0(ssrms0_out[15]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[14]), .Y(n4185) );
  NOR2XLTS U5021 ( .A(n4243), .B(n4224), .Y(n4184) );
  AO22XLTS U5022 ( .A0(n4293), .A1(aluone_out[14]), .B0(n4227), .B1(n4179), 
        .Y(n4180) );
  AOI211XLTS U5023 ( .A0(ssrms0_out[13]), .A1(n4274), .B0(n4297), .C0(n4180), 
        .Y(n4183) );
  INVX2TS U5024 ( .A(n4184), .Y(n4181) );
  AOI32X1TS U5025 ( .A0(n4185), .A1(n4184), .A2(n4183), .B0(n4182), .B1(n4181), 
        .Y(n1893) );
  AOI22X1TS U5026 ( .A0(ssrms0_out[14]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[13]), .Y(n4192) );
  NOR2XLTS U5027 ( .A(n4252), .B(n4224), .Y(n4191) );
  AO22XLTS U5028 ( .A0(n4293), .A1(aluone_out[13]), .B0(n4227), .B1(n4186), 
        .Y(n4187) );
  AOI211XLTS U5029 ( .A0(ssrms0_out[12]), .A1(n4274), .B0(n4297), .C0(n4187), 
        .Y(n4190) );
  INVX2TS U5030 ( .A(n4191), .Y(n4188) );
  AOI32X1TS U5031 ( .A0(n4192), .A1(n4191), .A2(n4190), .B0(n4189), .B1(n4188), 
        .Y(n1892) );
  AOI22X1TS U5032 ( .A0(ssrms0_out[11]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[12]), .Y(n4199) );
  NOR2XLTS U5033 ( .A(n4261), .B(n4224), .Y(n4198) );
  AO22XLTS U5034 ( .A0(n4293), .A1(aluone_out[12]), .B0(n4227), .B1(n4193), 
        .Y(n4194) );
  AOI211XLTS U5035 ( .A0(ssrms0_out[13]), .A1(n4298), .B0(n4297), .C0(n4194), 
        .Y(n4197) );
  INVX2TS U5036 ( .A(n4198), .Y(n4195) );
  AOI32X1TS U5037 ( .A0(n4199), .A1(n4198), .A2(n4197), .B0(n4196), .B1(n4195), 
        .Y(n1891) );
  AOI22X1TS U5038 ( .A0(ssrms0_out[10]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[11]), .Y(n4207) );
  NOR2XLTS U5039 ( .A(n4270), .B(n4224), .Y(n4206) );
  OAI22X1TS U5040 ( .A0(n4201), .A1(n4282), .B0(n4209), .B1(n4200), .Y(n4202)
         );
  AOI211XLTS U5041 ( .A0(ssrms0_out[12]), .A1(n4298), .B0(n4297), .C0(n4202), 
        .Y(n4205) );
  INVX2TS U5042 ( .A(n4206), .Y(n4203) );
  AOI32X1TS U5043 ( .A0(n4207), .A1(n4206), .A2(n4205), .B0(n4204), .B1(n4203), 
        .Y(n1890) );
  AOI22X1TS U5044 ( .A0(ssrms0_out[11]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[10]), .Y(n4216) );
  NOR2XLTS U5045 ( .A(n4280), .B(n4224), .Y(n4215) );
  OAI22X1TS U5046 ( .A0(n4210), .A1(n4282), .B0(n4209), .B1(n4208), .Y(n4211)
         );
  AOI211XLTS U5047 ( .A0(ssrms0_out[9]), .A1(n4274), .B0(n4297), .C0(n4211), 
        .Y(n4214) );
  INVX2TS U5048 ( .A(n4215), .Y(n4212) );
  AOI32X1TS U5049 ( .A0(n4216), .A1(n4215), .A2(n4214), .B0(n4213), .B1(n4212), 
        .Y(n1889) );
  AOI22X1TS U5050 ( .A0(ssrms0_out[8]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[9]), .Y(n4223) );
  NOR2XLTS U5051 ( .A(n4292), .B(n4224), .Y(n4222) );
  AO22XLTS U5052 ( .A0(n4293), .A1(aluone_out[9]), .B0(n4227), .B1(n4217), .Y(
        n4218) );
  AOI211XLTS U5053 ( .A0(ssrms0_out[10]), .A1(n4298), .B0(n4297), .C0(n4218), 
        .Y(n4221) );
  INVX2TS U5054 ( .A(n4222), .Y(n4219) );
  AOI32X1TS U5055 ( .A0(n4223), .A1(n4222), .A2(n4221), .B0(n4220), .B1(n4219), 
        .Y(n1888) );
  AOI22X1TS U5056 ( .A0(ssrms0_out[7]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[8]), .Y(n4233) );
  NOR2XLTS U5057 ( .A(n4225), .B(n4224), .Y(n4232) );
  AO22XLTS U5058 ( .A0(n4227), .A1(n4226), .B0(n4293), .B1(aluone_out[8]), .Y(
        n4228) );
  AOI211XLTS U5059 ( .A0(ssrms0_out[9]), .A1(n4298), .B0(n4297), .C0(n4228), 
        .Y(n4231) );
  INVX2TS U5060 ( .A(ssrms0_out[8]), .Y(n4230) );
  INVX2TS U5061 ( .A(n4232), .Y(n4229) );
  AOI32X1TS U5062 ( .A0(n4233), .A1(n4232), .A2(n4231), .B0(n4230), .B1(n4229), 
        .Y(n1887) );
  AOI22X1TS U5063 ( .A0(ssrms0_out[8]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[7]), .Y(n4242) );
  NOR2XLTS U5064 ( .A(n4234), .B(n4291), .Y(n4241) );
  OAI22X1TS U5065 ( .A0(n4236), .A1(n4282), .B0(n4235), .B1(n4294), .Y(n4237)
         );
  AOI211XLTS U5066 ( .A0(ssrms0_out[6]), .A1(n4274), .B0(n4297), .C0(n4237), 
        .Y(n4240) );
  INVX2TS U5067 ( .A(n4241), .Y(n4238) );
  AOI32X1TS U5068 ( .A0(n4242), .A1(n4241), .A2(n4240), .B0(n4239), .B1(n4238), 
        .Y(n1886) );
  AOI22X1TS U5069 ( .A0(ssrms0_out[5]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[6]), .Y(n4251) );
  NOR2XLTS U5070 ( .A(n4243), .B(n4291), .Y(n4250) );
  OAI22X1TS U5071 ( .A0(n4245), .A1(n4294), .B0(n4244), .B1(n4282), .Y(n4246)
         );
  AOI211XLTS U5072 ( .A0(ssrms0_out[7]), .A1(n4298), .B0(n4297), .C0(n4246), 
        .Y(n4249) );
  INVX2TS U5073 ( .A(n4250), .Y(n4247) );
  AOI32X1TS U5074 ( .A0(n4251), .A1(n4250), .A2(n4249), .B0(n4248), .B1(n4247), 
        .Y(n1885) );
  AOI22X1TS U5075 ( .A0(ssrms0_out[4]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[5]), .Y(n4260) );
  NOR2XLTS U5076 ( .A(n4252), .B(n4291), .Y(n4259) );
  OAI22X1TS U5077 ( .A0(n4254), .A1(n4294), .B0(n4253), .B1(n4282), .Y(n4255)
         );
  AOI211XLTS U5078 ( .A0(ssrms0_out[6]), .A1(n4298), .B0(n4297), .C0(n4255), 
        .Y(n4258) );
  INVX2TS U5079 ( .A(n4259), .Y(n4256) );
  AOI32X1TS U5080 ( .A0(n4260), .A1(n4259), .A2(n4258), .B0(n4257), .B1(n4256), 
        .Y(n1884) );
  AOI22X1TS U5081 ( .A0(ssrms0_out[5]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[4]), .Y(n4269) );
  NOR2XLTS U5082 ( .A(n4261), .B(n4291), .Y(n4268) );
  OAI22X1TS U5083 ( .A0(n4263), .A1(n4294), .B0(n4262), .B1(n4282), .Y(n4264)
         );
  AOI211XLTS U5084 ( .A0(ssrms0_out[3]), .A1(n4274), .B0(n4297), .C0(n4264), 
        .Y(n4267) );
  INVX2TS U5085 ( .A(n4268), .Y(n4265) );
  AOI32X1TS U5086 ( .A0(n4269), .A1(n4268), .A2(n4267), .B0(n4266), .B1(n4265), 
        .Y(n1883) );
  AOI22X1TS U5087 ( .A0(ssrms0_out[4]), .A1(n4298), .B0(n4290), .B1(
        mult1_out[3]), .Y(n4279) );
  NOR2XLTS U5088 ( .A(n4270), .B(n4291), .Y(n4278) );
  AO22XLTS U5089 ( .A0(n4293), .A1(aluone_out[3]), .B0(n4272), .B1(n4271), .Y(
        n4273) );
  AOI211XLTS U5090 ( .A0(ssrms0_out[2]), .A1(n4274), .B0(n4297), .C0(n4273), 
        .Y(n4277) );
  INVX2TS U5091 ( .A(n4278), .Y(n4275) );
  AOI32X1TS U5092 ( .A0(n4279), .A1(n4278), .A2(n4277), .B0(n4276), .B1(n4275), 
        .Y(n1882) );
  AOI22X1TS U5093 ( .A0(ssrms0_out[1]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[2]), .Y(n4289) );
  NOR2XLTS U5094 ( .A(n4280), .B(n4291), .Y(n4288) );
  OAI22X1TS U5095 ( .A0(n4283), .A1(n4282), .B0(n4281), .B1(n4294), .Y(n4284)
         );
  AOI211XLTS U5096 ( .A0(ssrms0_out[3]), .A1(n4298), .B0(n4297), .C0(n4284), 
        .Y(n4287) );
  INVX2TS U5097 ( .A(n4288), .Y(n4285) );
  AOI32X1TS U5098 ( .A0(n4289), .A1(n4288), .A2(n4287), .B0(n4286), .B1(n4285), 
        .Y(n1881) );
  AOI22X1TS U5099 ( .A0(ssrms0_out[0]), .A1(n4274), .B0(n4290), .B1(
        mult1_out[1]), .Y(n4303) );
  NOR2XLTS U5100 ( .A(n4292), .B(n4291), .Y(n4302) );
  OAI2BB2XLTS U5101 ( .B0(n4295), .B1(n4294), .A0N(aluone_out[1]), .A1N(n4293), 
        .Y(n4296) );
  AOI211XLTS U5102 ( .A0(ssrms0_out[2]), .A1(n4298), .B0(n4297), .C0(n4296), 
        .Y(n4301) );
  INVX2TS U5103 ( .A(n4302), .Y(n4299) );
  AOI32X1TS U5104 ( .A0(n4303), .A1(n4302), .A2(n4301), .B0(n4300), .B1(n4299), 
        .Y(n1880) );
  AOI22X1TS U5105 ( .A0(n1985), .A1(srmp_out[63]), .B0(n4407), .B1(
        srmp_out[62]), .Y(n4306) );
  NAND2X1TS U5106 ( .A(n4306), .B(n4305), .Y(n1878) );
  AOI22X1TS U5107 ( .A0(n4413), .A1(mult2_out[53]), .B0(n1985), .B1(
        srmp_out[53]), .Y(n4308) );
  AOI22X1TS U5108 ( .A0(n4407), .A1(srmp_out[52]), .B0(n4412), .B1(
        srmp_out[54]), .Y(n4307) );
  NAND2X1TS U5109 ( .A(n4308), .B(n4307), .Y(n1868) );
  AOI22X1TS U5110 ( .A0(n1985), .A1(srmp_out[52]), .B0(n4407), .B1(
        srmp_out[51]), .Y(n4310) );
  AOI22X1TS U5111 ( .A0(n4413), .A1(mult2_out[52]), .B0(n4412), .B1(
        srmp_out[53]), .Y(n4309) );
  NAND2X1TS U5112 ( .A(n4310), .B(n4309), .Y(n1867) );
  AOI22X1TS U5113 ( .A0(n1985), .A1(srmp_out[51]), .B0(n4407), .B1(
        srmp_out[50]), .Y(n4312) );
  AOI22X1TS U5114 ( .A0(n4413), .A1(mult2_out[51]), .B0(n4412), .B1(
        srmp_out[52]), .Y(n4311) );
  NAND2X1TS U5115 ( .A(n4312), .B(n4311), .Y(n1866) );
  AOI22X1TS U5116 ( .A0(n1985), .A1(srmp_out[50]), .B0(n4412), .B1(
        srmp_out[51]), .Y(n4314) );
  AOI22X1TS U5117 ( .A0(n4413), .A1(mult2_out[50]), .B0(n4407), .B1(
        srmp_out[49]), .Y(n4313) );
  NAND2X1TS U5118 ( .A(n4314), .B(n4313), .Y(n1865) );
  AOI22X1TS U5119 ( .A0(n4407), .A1(srmp_out[48]), .B0(n4412), .B1(
        srmp_out[50]), .Y(n4316) );
  AOI22X1TS U5120 ( .A0(n4413), .A1(mult2_out[49]), .B0(n1985), .B1(
        srmp_out[49]), .Y(n4315) );
  NAND2X1TS U5121 ( .A(n4316), .B(n4315), .Y(n1864) );
  AOI22X1TS U5122 ( .A0(n4413), .A1(mult2_out[48]), .B0(n4407), .B1(
        srmp_out[47]), .Y(n4318) );
  AOI22X1TS U5123 ( .A0(n1985), .A1(srmp_out[48]), .B0(n4412), .B1(
        srmp_out[49]), .Y(n4317) );
  NAND2X1TS U5124 ( .A(n4318), .B(n4317), .Y(n1863) );
  AOI22X1TS U5125 ( .A0(n4413), .A1(mult2_out[47]), .B0(n4407), .B1(
        srmp_out[46]), .Y(n4320) );
  AOI22X1TS U5126 ( .A0(n1985), .A1(srmp_out[47]), .B0(n4412), .B1(
        srmp_out[48]), .Y(n4319) );
  NAND2X1TS U5127 ( .A(n4320), .B(n4319), .Y(n1862) );
  AOI22X1TS U5128 ( .A0(n4407), .A1(srmp_out[45]), .B0(n4412), .B1(
        srmp_out[47]), .Y(n4322) );
  AOI22X1TS U5129 ( .A0(n4413), .A1(mult2_out[46]), .B0(n1985), .B1(
        srmp_out[46]), .Y(n4321) );
  NAND2X1TS U5130 ( .A(n4322), .B(n4321), .Y(n1861) );
  AOI22X1TS U5131 ( .A0(n1985), .A1(srmp_out[45]), .B0(n4412), .B1(
        srmp_out[46]), .Y(n4324) );
  AOI22X1TS U5132 ( .A0(n4413), .A1(mult2_out[45]), .B0(n4407), .B1(
        srmp_out[44]), .Y(n4323) );
  NAND2X1TS U5133 ( .A(n4324), .B(n4323), .Y(n1860) );
  AOI22X1TS U5134 ( .A0(n4407), .A1(srmp_out[43]), .B0(n4412), .B1(
        srmp_out[45]), .Y(n4326) );
  AOI22X1TS U5135 ( .A0(n4413), .A1(mult2_out[44]), .B0(n1985), .B1(
        srmp_out[44]), .Y(n4325) );
  NAND2X1TS U5136 ( .A(n4326), .B(n4325), .Y(n1859) );
  AOI22X1TS U5137 ( .A0(n4413), .A1(mult2_out[43]), .B0(n1985), .B1(
        srmp_out[43]), .Y(n4328) );
  AOI22X1TS U5138 ( .A0(n4407), .A1(srmp_out[42]), .B0(n4412), .B1(
        srmp_out[44]), .Y(n4327) );
  NAND2X1TS U5139 ( .A(n4328), .B(n4327), .Y(n1858) );
  AOI22X1TS U5140 ( .A0(n1985), .A1(srmp_out[42]), .B0(n4407), .B1(
        srmp_out[41]), .Y(n4330) );
  AOI22X1TS U5141 ( .A0(n4413), .A1(mult2_out[42]), .B0(n4412), .B1(
        srmp_out[43]), .Y(n4329) );
  NAND2X1TS U5142 ( .A(n4330), .B(n4329), .Y(n1857) );
  AOI22X1TS U5143 ( .A0(n4413), .A1(mult2_out[41]), .B0(n4412), .B1(
        srmp_out[42]), .Y(n4332) );
  AOI22X1TS U5144 ( .A0(n1985), .A1(srmp_out[41]), .B0(n4407), .B1(
        srmp_out[40]), .Y(n4331) );
  NAND2X1TS U5145 ( .A(n4332), .B(n4331), .Y(n1856) );
  AOI22X1TS U5146 ( .A0(n1985), .A1(srmp_out[40]), .B0(n4407), .B1(
        srmp_out[39]), .Y(n4334) );
  AOI22X1TS U5147 ( .A0(n4413), .A1(mult2_out[40]), .B0(n4412), .B1(
        srmp_out[41]), .Y(n4333) );
  NAND2X1TS U5148 ( .A(n4334), .B(n4333), .Y(n1855) );
  AOI22X1TS U5149 ( .A0(n4413), .A1(mult2_out[39]), .B0(n1985), .B1(
        srmp_out[39]), .Y(n4336) );
  AOI22X1TS U5150 ( .A0(n4407), .A1(srmp_out[38]), .B0(n4412), .B1(
        srmp_out[40]), .Y(n4335) );
  NAND2X1TS U5151 ( .A(n4336), .B(n4335), .Y(n1854) );
  AOI22X1TS U5152 ( .A0(n4407), .A1(srmp_out[37]), .B0(n4412), .B1(
        srmp_out[39]), .Y(n4338) );
  AOI22X1TS U5153 ( .A0(n4413), .A1(mult2_out[38]), .B0(n1985), .B1(
        srmp_out[38]), .Y(n4337) );
  NAND2X1TS U5154 ( .A(n4338), .B(n4337), .Y(n1853) );
  AOI22X1TS U5155 ( .A0(n4413), .A1(mult2_out[37]), .B0(n4407), .B1(
        srmp_out[36]), .Y(n4340) );
  AOI22X1TS U5156 ( .A0(n1985), .A1(srmp_out[37]), .B0(n4412), .B1(
        srmp_out[38]), .Y(n4339) );
  NAND2X1TS U5157 ( .A(n4340), .B(n4339), .Y(n1852) );
  AOI22X1TS U5158 ( .A0(n4413), .A1(mult2_out[36]), .B0(n4412), .B1(
        srmp_out[37]), .Y(n4342) );
  AOI22X1TS U5159 ( .A0(n1985), .A1(srmp_out[36]), .B0(n4407), .B1(
        srmp_out[35]), .Y(n4341) );
  NAND2X1TS U5160 ( .A(n4342), .B(n4341), .Y(n1851) );
  AOI22X1TS U5161 ( .A0(n4413), .A1(mult2_out[35]), .B0(n4407), .B1(
        srmp_out[34]), .Y(n4344) );
  AOI22X1TS U5162 ( .A0(n1985), .A1(srmp_out[35]), .B0(n4412), .B1(
        srmp_out[36]), .Y(n4343) );
  NAND2X1TS U5163 ( .A(n4344), .B(n4343), .Y(n1850) );
  AOI22X1TS U5164 ( .A0(n4413), .A1(mult2_out[34]), .B0(n4407), .B1(
        srmp_out[33]), .Y(n4346) );
  AOI22X1TS U5165 ( .A0(n1985), .A1(srmp_out[34]), .B0(n4412), .B1(
        srmp_out[35]), .Y(n4345) );
  NAND2X1TS U5166 ( .A(n4346), .B(n4345), .Y(n1849) );
  AOI22X1TS U5167 ( .A0(n4413), .A1(mult2_out[33]), .B0(n1985), .B1(
        srmp_out[33]), .Y(n4348) );
  AOI22X1TS U5168 ( .A0(n4407), .A1(srmp_out[32]), .B0(n4412), .B1(
        srmp_out[34]), .Y(n4347) );
  NAND2X1TS U5169 ( .A(n4348), .B(n4347), .Y(n1848) );
  AOI22X1TS U5170 ( .A0(n1985), .A1(srmp_out[32]), .B0(n4407), .B1(
        srmp_out[31]), .Y(n4350) );
  AOI22X1TS U5171 ( .A0(n4413), .A1(mult2_out[32]), .B0(n4412), .B1(
        srmp_out[33]), .Y(n4349) );
  NAND2X1TS U5172 ( .A(n4350), .B(n4349), .Y(n1847) );
  AOI22X1TS U5173 ( .A0(n4413), .A1(mult2_out[31]), .B0(n1985), .B1(
        srmp_out[31]), .Y(n4352) );
  AOI22X1TS U5174 ( .A0(n4407), .A1(srmp_out[30]), .B0(n4412), .B1(
        srmp_out[32]), .Y(n4351) );
  NAND2X1TS U5175 ( .A(n4352), .B(n4351), .Y(n1846) );
  AOI22X1TS U5176 ( .A0(n1985), .A1(srmp_out[30]), .B0(n4412), .B1(
        srmp_out[31]), .Y(n4354) );
  AOI22X1TS U5177 ( .A0(n4413), .A1(mult2_out[30]), .B0(n4407), .B1(
        srmp_out[29]), .Y(n4353) );
  NAND2X1TS U5178 ( .A(n4354), .B(n4353), .Y(n1845) );
  AOI22X1TS U5179 ( .A0(n1985), .A1(srmp_out[29]), .B0(n4412), .B1(
        srmp_out[30]), .Y(n4356) );
  AOI22X1TS U5180 ( .A0(n4413), .A1(mult2_out[29]), .B0(n4407), .B1(
        srmp_out[28]), .Y(n4355) );
  NAND2X1TS U5181 ( .A(n4356), .B(n4355), .Y(n1844) );
  AOI22X1TS U5182 ( .A0(n1985), .A1(srmp_out[28]), .B0(n4407), .B1(
        srmp_out[27]), .Y(n4358) );
  AOI22X1TS U5183 ( .A0(n4413), .A1(mult2_out[28]), .B0(n4412), .B1(
        srmp_out[29]), .Y(n4357) );
  NAND2X1TS U5184 ( .A(n4358), .B(n4357), .Y(n1843) );
  AOI22X1TS U5185 ( .A0(n4407), .A1(srmp_out[26]), .B0(n4412), .B1(
        srmp_out[28]), .Y(n4360) );
  AOI22X1TS U5186 ( .A0(n4413), .A1(mult2_out[27]), .B0(n1985), .B1(
        srmp_out[27]), .Y(n4359) );
  NAND2X1TS U5187 ( .A(n4360), .B(n4359), .Y(n1842) );
  AOI22X1TS U5188 ( .A0(n4413), .A1(mult2_out[26]), .B0(n4412), .B1(
        srmp_out[27]), .Y(n4362) );
  AOI22X1TS U5189 ( .A0(n1985), .A1(srmp_out[26]), .B0(n4407), .B1(
        srmp_out[25]), .Y(n4361) );
  NAND2X1TS U5190 ( .A(n4362), .B(n4361), .Y(n1841) );
  AOI22X1TS U5191 ( .A0(n1985), .A1(srmp_out[25]), .B0(n4407), .B1(
        srmp_out[24]), .Y(n4364) );
  AOI22X1TS U5192 ( .A0(n4413), .A1(mult2_out[25]), .B0(n4412), .B1(
        srmp_out[26]), .Y(n4363) );
  NAND2X1TS U5193 ( .A(n4364), .B(n4363), .Y(n1840) );
  AOI22X1TS U5194 ( .A0(n4413), .A1(mult2_out[24]), .B0(n1985), .B1(
        srmp_out[24]), .Y(n4366) );
  AOI22X1TS U5195 ( .A0(n4407), .A1(srmp_out[23]), .B0(n4412), .B1(
        srmp_out[25]), .Y(n4365) );
  NAND2X1TS U5196 ( .A(n4366), .B(n4365), .Y(n1839) );
  AOI22X1TS U5197 ( .A0(n4413), .A1(mult2_out[23]), .B0(n1985), .B1(
        srmp_out[23]), .Y(n4368) );
  AOI22X1TS U5198 ( .A0(n4407), .A1(srmp_out[22]), .B0(n4412), .B1(
        srmp_out[24]), .Y(n4367) );
  NAND2X1TS U5199 ( .A(n4368), .B(n4367), .Y(n1838) );
  AOI22X1TS U5200 ( .A0(n4407), .A1(srmp_out[21]), .B0(n4412), .B1(
        srmp_out[23]), .Y(n4370) );
  AOI22X1TS U5201 ( .A0(n4413), .A1(mult2_out[22]), .B0(n1985), .B1(
        srmp_out[22]), .Y(n4369) );
  NAND2X1TS U5202 ( .A(n4370), .B(n4369), .Y(n1837) );
  AOI22X1TS U5203 ( .A0(n4413), .A1(mult2_out[21]), .B0(n1985), .B1(
        srmp_out[21]), .Y(n4372) );
  AOI22X1TS U5204 ( .A0(n4407), .A1(srmp_out[20]), .B0(n4412), .B1(
        srmp_out[22]), .Y(n4371) );
  NAND2X1TS U5205 ( .A(n4372), .B(n4371), .Y(n1836) );
  AOI22X1TS U5206 ( .A0(n4407), .A1(srmp_out[19]), .B0(n4412), .B1(
        srmp_out[21]), .Y(n4374) );
  AOI22X1TS U5207 ( .A0(n4413), .A1(mult2_out[20]), .B0(n1985), .B1(
        srmp_out[20]), .Y(n4373) );
  NAND2X1TS U5208 ( .A(n4374), .B(n4373), .Y(n1835) );
  AOI22X1TS U5209 ( .A0(n4407), .A1(srmp_out[18]), .B0(n4412), .B1(
        srmp_out[20]), .Y(n4376) );
  AOI22X1TS U5210 ( .A0(n4413), .A1(mult2_out[19]), .B0(n1985), .B1(
        srmp_out[19]), .Y(n4375) );
  NAND2X1TS U5211 ( .A(n4376), .B(n4375), .Y(n1834) );
  AOI22X1TS U5212 ( .A0(n4413), .A1(mult2_out[18]), .B0(n4412), .B1(
        srmp_out[19]), .Y(n4378) );
  AOI22X1TS U5213 ( .A0(n1985), .A1(srmp_out[18]), .B0(n4407), .B1(
        srmp_out[17]), .Y(n4377) );
  NAND2X1TS U5214 ( .A(n4378), .B(n4377), .Y(n1833) );
  AOI22X1TS U5215 ( .A0(n4413), .A1(mult2_out[17]), .B0(n4407), .B1(
        srmp_out[16]), .Y(n4380) );
  AOI22X1TS U5216 ( .A0(n1985), .A1(srmp_out[17]), .B0(n4412), .B1(
        srmp_out[18]), .Y(n4379) );
  NAND2X1TS U5217 ( .A(n4380), .B(n4379), .Y(n1832) );
  AOI22X1TS U5218 ( .A0(n4413), .A1(mult2_out[16]), .B0(n4407), .B1(
        srmp_out[15]), .Y(n4382) );
  AOI22X1TS U5219 ( .A0(n1985), .A1(srmp_out[16]), .B0(n4412), .B1(
        srmp_out[17]), .Y(n4381) );
  NAND2X1TS U5220 ( .A(n4382), .B(n4381), .Y(n1831) );
  AOI22X1TS U5221 ( .A0(n1985), .A1(srmp_out[15]), .B0(n4412), .B1(
        srmp_out[16]), .Y(n4384) );
  AOI22X1TS U5222 ( .A0(n4413), .A1(mult2_out[15]), .B0(n4407), .B1(
        srmp_out[14]), .Y(n4383) );
  NAND2X1TS U5223 ( .A(n4384), .B(n4383), .Y(n1830) );
  AOI22X1TS U5224 ( .A0(n4413), .A1(mult2_out[14]), .B0(n4412), .B1(
        srmp_out[15]), .Y(n4386) );
  AOI22X1TS U5225 ( .A0(n1985), .A1(srmp_out[14]), .B0(n4407), .B1(
        srmp_out[13]), .Y(n4385) );
  NAND2X1TS U5226 ( .A(n4386), .B(n4385), .Y(n1829) );
  AOI22X1TS U5227 ( .A0(n1985), .A1(srmp_out[13]), .B0(n4412), .B1(
        srmp_out[14]), .Y(n4388) );
  AOI22X1TS U5228 ( .A0(n4413), .A1(mult2_out[13]), .B0(n4407), .B1(
        srmp_out[12]), .Y(n4387) );
  NAND2X1TS U5229 ( .A(n4388), .B(n4387), .Y(n1828) );
  AOI22X1TS U5230 ( .A0(n1985), .A1(srmp_out[12]), .B0(n4407), .B1(
        srmp_out[11]), .Y(n4390) );
  AOI22X1TS U5231 ( .A0(n4413), .A1(mult2_out[12]), .B0(n4412), .B1(
        srmp_out[13]), .Y(n4389) );
  NAND2X1TS U5232 ( .A(n4390), .B(n4389), .Y(n1827) );
  AOI22X1TS U5233 ( .A0(n1985), .A1(srmp_out[11]), .B0(n4407), .B1(
        srmp_out[10]), .Y(n4392) );
  AOI22X1TS U5234 ( .A0(n4413), .A1(mult2_out[11]), .B0(n4412), .B1(
        srmp_out[12]), .Y(n4391) );
  NAND2X1TS U5235 ( .A(n4392), .B(n4391), .Y(n1826) );
  AOI22X1TS U5236 ( .A0(n4413), .A1(mult2_out[10]), .B0(n4412), .B1(
        srmp_out[11]), .Y(n4394) );
  AOI22X1TS U5237 ( .A0(n1985), .A1(srmp_out[10]), .B0(n4407), .B1(srmp_out[9]), .Y(n4393) );
  NAND2X1TS U5238 ( .A(n4394), .B(n4393), .Y(n1825) );
  AOI22X1TS U5239 ( .A0(n4413), .A1(mult2_out[9]), .B0(n1985), .B1(srmp_out[9]), .Y(n4396) );
  AOI22X1TS U5240 ( .A0(n4407), .A1(srmp_out[8]), .B0(n4412), .B1(srmp_out[10]), .Y(n4395) );
  NAND2X1TS U5241 ( .A(n4396), .B(n4395), .Y(n1824) );
  AOI22X1TS U5242 ( .A0(n1985), .A1(srmp_out[8]), .B0(n4407), .B1(srmp_out[7]), 
        .Y(n4398) );
  AOI22X1TS U5243 ( .A0(n4413), .A1(mult2_out[8]), .B0(n4412), .B1(srmp_out[9]), .Y(n4397) );
  NAND2X1TS U5244 ( .A(n4398), .B(n4397), .Y(n1823) );
  AOI22X1TS U5245 ( .A0(n1985), .A1(srmp_out[7]), .B0(n4412), .B1(srmp_out[8]), 
        .Y(n4400) );
  AOI22X1TS U5246 ( .A0(n4413), .A1(mult2_out[7]), .B0(n4407), .B1(srmp_out[6]), .Y(n4399) );
  NAND2X1TS U5247 ( .A(n4400), .B(n4399), .Y(n1822) );
  AOI22X1TS U5248 ( .A0(n1985), .A1(srmp_out[6]), .B0(n4412), .B1(srmp_out[7]), 
        .Y(n4402) );
  AOI22X1TS U5249 ( .A0(n4413), .A1(mult2_out[6]), .B0(n4407), .B1(srmp_out[5]), .Y(n4401) );
  NAND2X1TS U5250 ( .A(n4402), .B(n4401), .Y(n1821) );
  AOI22X1TS U5251 ( .A0(n1985), .A1(srmp_out[5]), .B0(n4407), .B1(srmp_out[4]), 
        .Y(n4404) );
  AOI22X1TS U5252 ( .A0(n4413), .A1(mult2_out[5]), .B0(n4412), .B1(srmp_out[6]), .Y(n4403) );
  NAND2X1TS U5253 ( .A(n4404), .B(n4403), .Y(n1820) );
  AOI22X1TS U5254 ( .A0(n4407), .A1(srmp_out[3]), .B0(n4412), .B1(srmp_out[5]), 
        .Y(n4406) );
  AOI22X1TS U5255 ( .A0(n4413), .A1(mult2_out[4]), .B0(n1985), .B1(srmp_out[4]), .Y(n4405) );
  NAND2X1TS U5256 ( .A(n4406), .B(n4405), .Y(n1819) );
  AOI22X1TS U5257 ( .A0(n4407), .A1(srmp_out[2]), .B0(n4412), .B1(srmp_out[4]), 
        .Y(n4409) );
  AOI22X1TS U5258 ( .A0(n4413), .A1(mult2_out[3]), .B0(n1985), .B1(srmp_out[3]), .Y(n4408) );
  NAND2X1TS U5259 ( .A(n4409), .B(n4408), .Y(n1818) );
  AOI22X1TS U5260 ( .A0(n4413), .A1(mult2_out[2]), .B0(n4407), .B1(srmp_out[1]), .Y(n4411) );
  AOI22X1TS U5261 ( .A0(n1985), .A1(srmp_out[2]), .B0(n4412), .B1(srmp_out[3]), 
        .Y(n4410) );
  NAND2X1TS U5262 ( .A(n4411), .B(n4410), .Y(n1817) );
  AOI22X1TS U5263 ( .A0(n4407), .A1(srmp_out[0]), .B0(n4412), .B1(srmp_out[2]), 
        .Y(n4415) );
  AOI22X1TS U5264 ( .A0(n4413), .A1(mult2_out[1]), .B0(n1985), .B1(srmp_out[1]), .Y(n4414) );
  NAND2X1TS U5265 ( .A(n4415), .B(n4414), .Y(n1816) );
  INVX2TS U5266 ( .A(\sr_mt[0] ), .Y(n4417) );
  AOI22X1TS U5267 ( .A0(srmt_out[31]), .A1(n4483), .B0(n4473), .B1(m5_out[31]), 
        .Y(n4416) );
  OAI2BB1X1TS U5268 ( .A0N(srmt_out[30]), .A1N(n4476), .B0(n4416), .Y(n1814)
         );
  AOI22X1TS U5269 ( .A0(srmt_out[31]), .A1(n4479), .B0(srmt_out[29]), .B1(
        n4476), .Y(n4420) );
  AOI22X1TS U5270 ( .A0(srmt_out[30]), .A1(n4483), .B0(n4473), .B1(m5_out[30]), 
        .Y(n4419) );
  NAND2X1TS U5271 ( .A(n4420), .B(n4419), .Y(n1813) );
  AOI22X1TS U5272 ( .A0(srmt_out[28]), .A1(n4476), .B0(n4473), .B1(m5_out[29]), 
        .Y(n4422) );
  AOI22X1TS U5273 ( .A0(srmt_out[30]), .A1(n4479), .B0(srmt_out[29]), .B1(
        n4483), .Y(n4421) );
  NAND2X1TS U5274 ( .A(n4422), .B(n4421), .Y(n1812) );
  AOI22X1TS U5275 ( .A0(srmt_out[28]), .A1(n4483), .B0(srmt_out[27]), .B1(
        n4476), .Y(n4424) );
  AOI22X1TS U5276 ( .A0(srmt_out[29]), .A1(n4479), .B0(n4473), .B1(m5_out[28]), 
        .Y(n4423) );
  NAND2X1TS U5277 ( .A(n4424), .B(n4423), .Y(n1811) );
  AOI22X1TS U5278 ( .A0(srmt_out[28]), .A1(n4479), .B0(n4473), .B1(m5_out[27]), 
        .Y(n4426) );
  AOI22X1TS U5279 ( .A0(srmt_out[27]), .A1(n4483), .B0(srmt_out[26]), .B1(
        n4476), .Y(n4425) );
  NAND2X1TS U5280 ( .A(n4426), .B(n4425), .Y(n1810) );
  AOI22X1TS U5281 ( .A0(srmt_out[25]), .A1(n4476), .B0(n4473), .B1(m5_out[26]), 
        .Y(n4428) );
  AOI22X1TS U5282 ( .A0(srmt_out[27]), .A1(n4479), .B0(srmt_out[26]), .B1(
        n4483), .Y(n4427) );
  NAND2X1TS U5283 ( .A(n4428), .B(n4427), .Y(n1809) );
  AOI22X1TS U5284 ( .A0(srmt_out[26]), .A1(n4479), .B0(srmt_out[25]), .B1(
        n4483), .Y(n4430) );
  AOI22X1TS U5285 ( .A0(srmt_out[24]), .A1(n4476), .B0(n4473), .B1(m5_out[25]), 
        .Y(n4429) );
  NAND2X1TS U5286 ( .A(n4430), .B(n4429), .Y(n1808) );
  AOI22X1TS U5287 ( .A0(srmt_out[24]), .A1(n4483), .B0(srmt_out[23]), .B1(
        n4476), .Y(n4432) );
  AOI22X1TS U5288 ( .A0(srmt_out[25]), .A1(n4479), .B0(n4473), .B1(m5_out[24]), 
        .Y(n4431) );
  NAND2X1TS U5289 ( .A(n4432), .B(n4431), .Y(n1807) );
  AOI22X1TS U5290 ( .A0(srmt_out[24]), .A1(n4479), .B0(srmt_out[22]), .B1(
        n4476), .Y(n4434) );
  AOI22X1TS U5291 ( .A0(srmt_out[23]), .A1(n4483), .B0(n4473), .B1(m5_out[23]), 
        .Y(n4433) );
  NAND2X1TS U5292 ( .A(n4434), .B(n4433), .Y(n1806) );
  AOI22X1TS U5293 ( .A0(srmt_out[21]), .A1(n4476), .B0(n4473), .B1(m5_out[22]), 
        .Y(n4436) );
  AOI22X1TS U5294 ( .A0(srmt_out[23]), .A1(n4479), .B0(srmt_out[22]), .B1(
        n4483), .Y(n4435) );
  NAND2X1TS U5295 ( .A(n4436), .B(n4435), .Y(n1805) );
  AOI22X1TS U5296 ( .A0(srmt_out[22]), .A1(n4479), .B0(srmt_out[20]), .B1(
        n4476), .Y(n4438) );
  AOI22X1TS U5297 ( .A0(srmt_out[21]), .A1(n4483), .B0(n4473), .B1(m5_out[21]), 
        .Y(n4437) );
  NAND2X1TS U5298 ( .A(n4438), .B(n4437), .Y(n1804) );
  AOI22X1TS U5299 ( .A0(srmt_out[21]), .A1(n4479), .B0(n4473), .B1(m5_out[20]), 
        .Y(n4440) );
  AOI22X1TS U5300 ( .A0(srmt_out[20]), .A1(n4483), .B0(srmt_out[19]), .B1(
        n4476), .Y(n4439) );
  NAND2X1TS U5301 ( .A(n4440), .B(n4439), .Y(n1803) );
  AOI22X1TS U5302 ( .A0(srmt_out[18]), .A1(n4476), .B0(n4473), .B1(m5_out[19]), 
        .Y(n4442) );
  AOI22X1TS U5303 ( .A0(srmt_out[20]), .A1(n4479), .B0(srmt_out[19]), .B1(
        n4483), .Y(n4441) );
  NAND2X1TS U5304 ( .A(n4442), .B(n4441), .Y(n1802) );
  AOI22X1TS U5305 ( .A0(srmt_out[17]), .A1(n4476), .B0(n4473), .B1(m5_out[18]), 
        .Y(n4444) );
  AOI22X1TS U5306 ( .A0(srmt_out[19]), .A1(n4479), .B0(srmt_out[18]), .B1(
        n4483), .Y(n4443) );
  NAND2X1TS U5307 ( .A(n4444), .B(n4443), .Y(n1801) );
  AOI22X1TS U5308 ( .A0(srmt_out[16]), .A1(n4476), .B0(n4473), .B1(m5_out[17]), 
        .Y(n4446) );
  AOI22X1TS U5309 ( .A0(srmt_out[18]), .A1(n4479), .B0(srmt_out[17]), .B1(
        n4483), .Y(n4445) );
  NAND2X1TS U5310 ( .A(n4446), .B(n4445), .Y(n1800) );
  AOI22X1TS U5311 ( .A0(srmt_out[17]), .A1(n4479), .B0(srmt_out[16]), .B1(
        n4483), .Y(n4448) );
  AOI22X1TS U5312 ( .A0(srmt_out[15]), .A1(n4476), .B0(n4473), .B1(m5_out[16]), 
        .Y(n4447) );
  NAND2X1TS U5313 ( .A(n4448), .B(n4447), .Y(n1799) );
  AOI22X1TS U5314 ( .A0(srmt_out[16]), .A1(n4479), .B0(srmt_out[15]), .B1(
        n4483), .Y(n4450) );
  AOI22X1TS U5315 ( .A0(srmt_out[14]), .A1(n4476), .B0(n4473), .B1(m5_out[15]), 
        .Y(n4449) );
  NAND2X1TS U5316 ( .A(n4450), .B(n4449), .Y(n1798) );
  AOI22X1TS U5317 ( .A0(srmt_out[15]), .A1(n4479), .B0(n4473), .B1(m5_out[14]), 
        .Y(n4452) );
  AOI22X1TS U5318 ( .A0(srmt_out[14]), .A1(n4483), .B0(srmt_out[13]), .B1(
        n4476), .Y(n4451) );
  NAND2X1TS U5319 ( .A(n4452), .B(n4451), .Y(n1797) );
  AOI22X1TS U5320 ( .A0(srmt_out[14]), .A1(n4479), .B0(srmt_out[12]), .B1(
        n4476), .Y(n4454) );
  AOI22X1TS U5321 ( .A0(srmt_out[13]), .A1(n4483), .B0(n4473), .B1(m5_out[13]), 
        .Y(n4453) );
  NAND2X1TS U5322 ( .A(n4454), .B(n4453), .Y(n1796) );
  AOI22X1TS U5323 ( .A0(srmt_out[13]), .A1(n4479), .B0(srmt_out[12]), .B1(
        n4483), .Y(n4456) );
  AOI22X1TS U5324 ( .A0(srmt_out[11]), .A1(n4476), .B0(n4473), .B1(m5_out[12]), 
        .Y(n4455) );
  NAND2X1TS U5325 ( .A(n4456), .B(n4455), .Y(n1795) );
  AOI22X1TS U5326 ( .A0(srmt_out[12]), .A1(n4479), .B0(srmt_out[11]), .B1(
        n4483), .Y(n4458) );
  AOI22X1TS U5327 ( .A0(srmt_out[10]), .A1(n4476), .B0(n4473), .B1(m5_out[11]), 
        .Y(n4457) );
  NAND2X1TS U5328 ( .A(n4458), .B(n4457), .Y(n1794) );
  AOI22X1TS U5329 ( .A0(srmt_out[10]), .A1(n4483), .B0(srmt_out[9]), .B1(n4476), .Y(n4460) );
  AOI22X1TS U5330 ( .A0(srmt_out[11]), .A1(n4479), .B0(n4473), .B1(m5_out[10]), 
        .Y(n4459) );
  NAND2X1TS U5331 ( .A(n4460), .B(n4459), .Y(n1793) );
  AOI22X1TS U5332 ( .A0(srmt_out[10]), .A1(n4479), .B0(srmt_out[8]), .B1(n4476), .Y(n4462) );
  AOI22X1TS U5333 ( .A0(srmt_out[9]), .A1(n4483), .B0(n4473), .B1(m5_out[9]), 
        .Y(n4461) );
  NAND2X1TS U5334 ( .A(n4462), .B(n4461), .Y(n1792) );
  AOI22X1TS U5335 ( .A0(srmt_out[9]), .A1(n4479), .B0(n4473), .B1(m5_out[8]), 
        .Y(n4464) );
  AOI22X1TS U5336 ( .A0(srmt_out[8]), .A1(n4483), .B0(srmt_out[7]), .B1(n4476), 
        .Y(n4463) );
  NAND2X1TS U5337 ( .A(n4464), .B(n4463), .Y(n1791) );
  AOI22X1TS U5338 ( .A0(srmt_out[8]), .A1(n4479), .B0(srmt_out[6]), .B1(n4476), 
        .Y(n4466) );
  AOI22X1TS U5339 ( .A0(srmt_out[7]), .A1(n4483), .B0(n4473), .B1(m5_out[7]), 
        .Y(n4465) );
  NAND2X1TS U5340 ( .A(n4466), .B(n4465), .Y(n1790) );
  AOI22X1TS U5341 ( .A0(srmt_out[6]), .A1(n4483), .B0(srmt_out[5]), .B1(n4476), 
        .Y(n4468) );
  AOI22X1TS U5342 ( .A0(srmt_out[7]), .A1(n4479), .B0(n4473), .B1(m5_out[6]), 
        .Y(n4467) );
  NAND2X1TS U5343 ( .A(n4468), .B(n4467), .Y(n1789) );
  AOI22X1TS U5344 ( .A0(srmt_out[5]), .A1(n4483), .B0(srmt_out[4]), .B1(n4476), 
        .Y(n4470) );
  AOI22X1TS U5345 ( .A0(srmt_out[6]), .A1(n4479), .B0(n4473), .B1(m5_out[5]), 
        .Y(n4469) );
  NAND2X1TS U5346 ( .A(n4470), .B(n4469), .Y(n1788) );
  AOI22X1TS U5347 ( .A0(srmt_out[5]), .A1(n4479), .B0(srmt_out[3]), .B1(n4476), 
        .Y(n4472) );
  AOI22X1TS U5348 ( .A0(srmt_out[4]), .A1(n4483), .B0(n4473), .B1(m5_out[4]), 
        .Y(n4471) );
  NAND2X1TS U5349 ( .A(n4472), .B(n4471), .Y(n1787) );
  AOI22X1TS U5350 ( .A0(srmt_out[3]), .A1(n4483), .B0(srmt_out[2]), .B1(n4476), 
        .Y(n4475) );
  AOI22X1TS U5351 ( .A0(srmt_out[4]), .A1(n4479), .B0(n4473), .B1(m5_out[3]), 
        .Y(n4474) );
  NAND2X1TS U5352 ( .A(n4475), .B(n4474), .Y(n1786) );
  AOI22X1TS U5353 ( .A0(srmt_out[2]), .A1(n4483), .B0(n4473), .B1(m5_out[2]), 
        .Y(n4478) );
  AOI22X1TS U5354 ( .A0(srmt_out[3]), .A1(n4479), .B0(srmt_out[1]), .B1(n4476), 
        .Y(n4477) );
  NAND2X1TS U5355 ( .A(n4478), .B(n4477), .Y(n1785) );
  AOI22X1TS U5356 ( .A0(srmt_out[1]), .A1(n4483), .B0(srmt_out[0]), .B1(n4476), 
        .Y(n4481) );
  AOI22X1TS U5357 ( .A0(srmt_out[2]), .A1(n4479), .B0(n4473), .B1(m5_out[1]), 
        .Y(n4480) );
  NAND2X1TS U5358 ( .A(n4481), .B(n4480), .Y(n1784) );
  AOI22X1TS U5359 ( .A0(srmt_out[1]), .A1(n4479), .B0(n4473), .B1(m5_out[0]), 
        .Y(n4482) );
  OAI2BB1X1TS U5360 ( .A0N(srmt_out[0]), .A1N(n4483), .B0(n4482), .Y(n1783) );
  AOI22X1TS U5361 ( .A0(n1987), .A1(srmq_out[63]), .B0(n4592), .B1(
        srmq_out[62]), .Y(n4486) );
  NAND2X1TS U5362 ( .A(n4486), .B(n4485), .Y(n1782) );
  AOI22X1TS U5363 ( .A0(mult2_out[53]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[52]), .Y(n4488) );
  AOI22X1TS U5364 ( .A0(n1987), .A1(srmq_out[53]), .B0(n4597), .B1(
        srmq_out[54]), .Y(n4487) );
  NAND2X1TS U5365 ( .A(n4488), .B(n4487), .Y(n1772) );
  AOI22X1TS U5366 ( .A0(n1987), .A1(srmq_out[52]), .B0(n4597), .B1(
        srmq_out[53]), .Y(n4490) );
  AOI22X1TS U5367 ( .A0(mult2_out[52]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[51]), .Y(n4489) );
  NAND2X1TS U5368 ( .A(n4490), .B(n4489), .Y(n1771) );
  AOI22X1TS U5369 ( .A0(mult2_out[51]), .A1(n4515), .B0(n4597), .B1(
        srmq_out[52]), .Y(n4492) );
  AOI22X1TS U5370 ( .A0(n1987), .A1(srmq_out[51]), .B0(n4592), .B1(
        srmq_out[50]), .Y(n4491) );
  NAND2X1TS U5371 ( .A(n4492), .B(n4491), .Y(n1770) );
  AOI22X1TS U5372 ( .A0(n4592), .A1(srmq_out[49]), .B0(n4597), .B1(
        srmq_out[51]), .Y(n4494) );
  AOI22X1TS U5373 ( .A0(mult2_out[50]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[50]), .Y(n4493) );
  NAND2X1TS U5374 ( .A(n4494), .B(n4493), .Y(n1769) );
  AOI22X1TS U5375 ( .A0(n1987), .A1(srmq_out[49]), .B0(n4592), .B1(
        srmq_out[48]), .Y(n4496) );
  AOI22X1TS U5376 ( .A0(mult2_out[49]), .A1(n4515), .B0(n4597), .B1(
        srmq_out[50]), .Y(n4495) );
  NAND2X1TS U5377 ( .A(n4496), .B(n4495), .Y(n1768) );
  AOI22X1TS U5378 ( .A0(n1987), .A1(srmq_out[48]), .B0(n4597), .B1(
        srmq_out[49]), .Y(n4498) );
  AOI22X1TS U5379 ( .A0(mult2_out[48]), .A1(n4515), .B0(n4592), .B1(
        srmq_out[47]), .Y(n4497) );
  NAND2X1TS U5380 ( .A(n4498), .B(n4497), .Y(n1767) );
  AOI22X1TS U5381 ( .A0(mult2_out[47]), .A1(n4515), .B0(n1987), .B1(
        srmq_out[47]), .Y(n4500) );
  AOI22X1TS U5382 ( .A0(n4592), .A1(srmq_out[46]), .B0(n4597), .B1(
        srmq_out[48]), .Y(n4499) );
  NAND2X1TS U5383 ( .A(n4500), .B(n4499), .Y(n1766) );
  AOI22X1TS U5384 ( .A0(n1987), .A1(srmq_out[46]), .B0(n4597), .B1(
        srmq_out[47]), .Y(n4502) );
  AOI22X1TS U5385 ( .A0(mult2_out[46]), .A1(n4515), .B0(n4592), .B1(
        srmq_out[45]), .Y(n4501) );
  NAND2X1TS U5386 ( .A(n4502), .B(n4501), .Y(n1765) );
  AOI22X1TS U5387 ( .A0(n4592), .A1(srmq_out[44]), .B0(n4597), .B1(
        srmq_out[46]), .Y(n4504) );
  AOI22X1TS U5388 ( .A0(mult2_out[45]), .A1(n4515), .B0(n1987), .B1(
        srmq_out[45]), .Y(n4503) );
  NAND2X1TS U5389 ( .A(n4504), .B(n4503), .Y(n1764) );
  AOI22X1TS U5390 ( .A0(n1987), .A1(srmq_out[44]), .B0(n4597), .B1(
        srmq_out[45]), .Y(n4506) );
  AOI22X1TS U5391 ( .A0(mult2_out[44]), .A1(n4515), .B0(n4592), .B1(
        srmq_out[43]), .Y(n4505) );
  NAND2X1TS U5392 ( .A(n4506), .B(n4505), .Y(n1763) );
  AOI22X1TS U5393 ( .A0(mult2_out[43]), .A1(n4515), .B0(n4592), .B1(
        srmq_out[42]), .Y(n4508) );
  AOI22X1TS U5394 ( .A0(n1987), .A1(srmq_out[43]), .B0(n4597), .B1(
        srmq_out[44]), .Y(n4507) );
  NAND2X1TS U5395 ( .A(n4508), .B(n4507), .Y(n1762) );
  AOI22X1TS U5396 ( .A0(mult2_out[42]), .A1(n4515), .B0(n1987), .B1(
        srmq_out[42]), .Y(n4510) );
  AOI22X1TS U5397 ( .A0(n4592), .A1(srmq_out[41]), .B0(n4597), .B1(
        srmq_out[43]), .Y(n4509) );
  NAND2X1TS U5398 ( .A(n4510), .B(n4509), .Y(n1761) );
  AOI22X1TS U5399 ( .A0(mult2_out[41]), .A1(n4515), .B0(n1987), .B1(
        srmq_out[41]), .Y(n4512) );
  AOI22X1TS U5400 ( .A0(n4592), .A1(srmq_out[40]), .B0(n4597), .B1(
        srmq_out[42]), .Y(n4511) );
  NAND2X1TS U5401 ( .A(n4512), .B(n4511), .Y(n1760) );
  AOI22X1TS U5402 ( .A0(n1987), .A1(srmq_out[40]), .B0(n4592), .B1(
        srmq_out[39]), .Y(n4514) );
  AOI22X1TS U5403 ( .A0(mult2_out[40]), .A1(n4515), .B0(n4597), .B1(
        srmq_out[41]), .Y(n4513) );
  NAND2X1TS U5404 ( .A(n4514), .B(n4513), .Y(n1759) );
  AOI22X1TS U5405 ( .A0(n1987), .A1(srmq_out[39]), .B0(n4597), .B1(
        srmq_out[40]), .Y(n4517) );
  AOI22X1TS U5406 ( .A0(mult2_out[39]), .A1(n4515), .B0(n4592), .B1(
        srmq_out[38]), .Y(n4516) );
  NAND2X1TS U5407 ( .A(n4517), .B(n4516), .Y(n1758) );
  AOI22X1TS U5408 ( .A0(mult2_out[38]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[38]), .Y(n4519) );
  AOI22X1TS U5409 ( .A0(n4592), .A1(srmq_out[37]), .B0(n4597), .B1(
        srmq_out[39]), .Y(n4518) );
  NAND2X1TS U5410 ( .A(n4519), .B(n4518), .Y(n1757) );
  AOI22X1TS U5411 ( .A0(n1987), .A1(srmq_out[37]), .B0(n4597), .B1(
        srmq_out[38]), .Y(n4521) );
  AOI22X1TS U5412 ( .A0(mult2_out[37]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[36]), .Y(n4520) );
  NAND2X1TS U5413 ( .A(n4521), .B(n4520), .Y(n1756) );
  AOI22X1TS U5414 ( .A0(mult2_out[36]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[35]), .Y(n4523) );
  AOI22X1TS U5415 ( .A0(n1987), .A1(srmq_out[36]), .B0(n4597), .B1(
        srmq_out[37]), .Y(n4522) );
  NAND2X1TS U5416 ( .A(n4523), .B(n4522), .Y(n1755) );
  AOI22X1TS U5417 ( .A0(mult2_out[35]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[34]), .Y(n4525) );
  AOI22X1TS U5418 ( .A0(n1987), .A1(srmq_out[35]), .B0(n4597), .B1(
        srmq_out[36]), .Y(n4524) );
  NAND2X1TS U5419 ( .A(n4525), .B(n4524), .Y(n1754) );
  AOI22X1TS U5420 ( .A0(n4592), .A1(srmq_out[33]), .B0(n4597), .B1(
        srmq_out[35]), .Y(n4527) );
  AOI22X1TS U5421 ( .A0(mult2_out[34]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[34]), .Y(n4526) );
  NAND2X1TS U5422 ( .A(n4527), .B(n4526), .Y(n1753) );
  AOI22X1TS U5423 ( .A0(n1987), .A1(srmq_out[33]), .B0(n4592), .B1(
        srmq_out[32]), .Y(n4529) );
  AOI22X1TS U5424 ( .A0(mult2_out[33]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[34]), .Y(n4528) );
  NAND2X1TS U5425 ( .A(n4529), .B(n4528), .Y(n1752) );
  AOI22X1TS U5426 ( .A0(n4592), .A1(srmq_out[31]), .B0(n4597), .B1(
        srmq_out[33]), .Y(n4531) );
  AOI22X1TS U5427 ( .A0(mult2_out[32]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[32]), .Y(n4530) );
  NAND2X1TS U5428 ( .A(n4531), .B(n4530), .Y(n1751) );
  AOI22X1TS U5429 ( .A0(n4592), .A1(srmq_out[30]), .B0(n4597), .B1(
        srmq_out[32]), .Y(n4533) );
  AOI22X1TS U5430 ( .A0(mult2_out[31]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[31]), .Y(n4532) );
  NAND2X1TS U5431 ( .A(n4533), .B(n4532), .Y(n1750) );
  AOI22X1TS U5432 ( .A0(mult2_out[30]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[31]), .Y(n4535) );
  AOI22X1TS U5433 ( .A0(n1987), .A1(srmq_out[30]), .B0(n4592), .B1(
        srmq_out[29]), .Y(n4534) );
  NAND2X1TS U5434 ( .A(n4535), .B(n4534), .Y(n1749) );
  AOI22X1TS U5435 ( .A0(mult2_out[29]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[29]), .Y(n4537) );
  AOI22X1TS U5436 ( .A0(n4592), .A1(srmq_out[28]), .B0(n4597), .B1(
        srmq_out[30]), .Y(n4536) );
  NAND2X1TS U5437 ( .A(n4537), .B(n4536), .Y(n1748) );
  AOI22X1TS U5438 ( .A0(n1987), .A1(srmq_out[28]), .B0(n4592), .B1(
        srmq_out[27]), .Y(n4539) );
  AOI22X1TS U5439 ( .A0(mult2_out[28]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[29]), .Y(n4538) );
  NAND2X1TS U5440 ( .A(n4539), .B(n4538), .Y(n1747) );
  AOI22X1TS U5441 ( .A0(n1987), .A1(srmq_out[27]), .B0(n4597), .B1(
        srmq_out[28]), .Y(n4541) );
  AOI22X1TS U5442 ( .A0(mult2_out[27]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[26]), .Y(n4540) );
  NAND2X1TS U5443 ( .A(n4541), .B(n4540), .Y(n1746) );
  AOI22X1TS U5444 ( .A0(mult2_out[26]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[27]), .Y(n4543) );
  AOI22X1TS U5445 ( .A0(n1987), .A1(srmq_out[26]), .B0(n4592), .B1(
        srmq_out[25]), .Y(n4542) );
  NAND2X1TS U5446 ( .A(n4543), .B(n4542), .Y(n1745) );
  AOI22X1TS U5447 ( .A0(mult2_out[25]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[25]), .Y(n4545) );
  AOI22X1TS U5448 ( .A0(n4592), .A1(srmq_out[24]), .B0(n4597), .B1(
        srmq_out[26]), .Y(n4544) );
  NAND2X1TS U5449 ( .A(n4545), .B(n4544), .Y(n1744) );
  AOI22X1TS U5450 ( .A0(mult2_out[24]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[25]), .Y(n4547) );
  AOI22X1TS U5451 ( .A0(n1987), .A1(srmq_out[24]), .B0(n4592), .B1(
        srmq_out[23]), .Y(n4546) );
  NAND2X1TS U5452 ( .A(n4547), .B(n4546), .Y(n1743) );
  AOI22X1TS U5453 ( .A0(mult2_out[23]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[23]), .Y(n4549) );
  AOI22X1TS U5454 ( .A0(n4592), .A1(srmq_out[22]), .B0(n4597), .B1(
        srmq_out[24]), .Y(n4548) );
  NAND2X1TS U5455 ( .A(n4549), .B(n4548), .Y(n1742) );
  AOI22X1TS U5456 ( .A0(n4592), .A1(srmq_out[21]), .B0(n4597), .B1(
        srmq_out[23]), .Y(n4551) );
  AOI22X1TS U5457 ( .A0(mult2_out[22]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[22]), .Y(n4550) );
  NAND2X1TS U5458 ( .A(n4551), .B(n4550), .Y(n1741) );
  AOI22X1TS U5459 ( .A0(n1987), .A1(srmq_out[21]), .B0(n4597), .B1(
        srmq_out[22]), .Y(n4553) );
  AOI22X1TS U5460 ( .A0(mult2_out[21]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[20]), .Y(n4552) );
  NAND2X1TS U5461 ( .A(n4553), .B(n4552), .Y(n1740) );
  AOI22X1TS U5462 ( .A0(mult2_out[20]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[19]), .Y(n4555) );
  AOI22X1TS U5463 ( .A0(n1987), .A1(srmq_out[20]), .B0(n4597), .B1(
        srmq_out[21]), .Y(n4554) );
  NAND2X1TS U5464 ( .A(n4555), .B(n4554), .Y(n1739) );
  AOI22X1TS U5465 ( .A0(mult2_out[19]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[19]), .Y(n4557) );
  AOI22X1TS U5466 ( .A0(n4592), .A1(srmq_out[18]), .B0(n4597), .B1(
        srmq_out[20]), .Y(n4556) );
  NAND2X1TS U5467 ( .A(n4557), .B(n4556), .Y(n1738) );
  AOI22X1TS U5468 ( .A0(mult2_out[18]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[18]), .Y(n4559) );
  AOI22X1TS U5469 ( .A0(n4592), .A1(srmq_out[17]), .B0(n4597), .B1(
        srmq_out[19]), .Y(n4558) );
  NAND2X1TS U5470 ( .A(n4559), .B(n4558), .Y(n1737) );
  AOI22X1TS U5471 ( .A0(n1987), .A1(srmq_out[17]), .B0(n4597), .B1(
        srmq_out[18]), .Y(n4561) );
  AOI22X1TS U5472 ( .A0(mult2_out[17]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[16]), .Y(n4560) );
  NAND2X1TS U5473 ( .A(n4561), .B(n4560), .Y(n1736) );
  AOI22X1TS U5474 ( .A0(mult2_out[16]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[15]), .Y(n4563) );
  AOI22X1TS U5475 ( .A0(n1987), .A1(srmq_out[16]), .B0(n4597), .B1(
        srmq_out[17]), .Y(n4562) );
  NAND2X1TS U5476 ( .A(n4563), .B(n4562), .Y(n1735) );
  AOI22X1TS U5477 ( .A0(n1987), .A1(srmq_out[15]), .B0(n4597), .B1(
        srmq_out[16]), .Y(n4565) );
  AOI22X1TS U5478 ( .A0(mult2_out[15]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[14]), .Y(n4564) );
  NAND2X1TS U5479 ( .A(n4565), .B(n4564), .Y(n1734) );
  AOI22X1TS U5480 ( .A0(n1987), .A1(srmq_out[14]), .B0(n4592), .B1(
        srmq_out[13]), .Y(n4567) );
  AOI22X1TS U5481 ( .A0(mult2_out[14]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[15]), .Y(n4566) );
  NAND2X1TS U5482 ( .A(n4567), .B(n4566), .Y(n1733) );
  AOI22X1TS U5483 ( .A0(mult2_out[13]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[13]), .Y(n4569) );
  AOI22X1TS U5484 ( .A0(n4592), .A1(srmq_out[12]), .B0(n4597), .B1(
        srmq_out[14]), .Y(n4568) );
  NAND2X1TS U5485 ( .A(n4569), .B(n4568), .Y(n1732) );
  AOI22X1TS U5486 ( .A0(n4592), .A1(srmq_out[11]), .B0(n4597), .B1(
        srmq_out[13]), .Y(n4571) );
  AOI22X1TS U5487 ( .A0(mult2_out[12]), .A1(n4595), .B0(n1987), .B1(
        srmq_out[12]), .Y(n4570) );
  NAND2X1TS U5488 ( .A(n4571), .B(n4570), .Y(n1731) );
  AOI22X1TS U5489 ( .A0(n1987), .A1(srmq_out[11]), .B0(n4597), .B1(
        srmq_out[12]), .Y(n4573) );
  AOI22X1TS U5490 ( .A0(mult2_out[11]), .A1(n4595), .B0(n4592), .B1(
        srmq_out[10]), .Y(n4572) );
  NAND2X1TS U5491 ( .A(n4573), .B(n4572), .Y(n1730) );
  AOI22X1TS U5492 ( .A0(mult2_out[10]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[11]), .Y(n4575) );
  AOI22X1TS U5493 ( .A0(n1987), .A1(srmq_out[10]), .B0(n4592), .B1(srmq_out[9]), .Y(n4574) );
  NAND2X1TS U5494 ( .A(n4575), .B(n4574), .Y(n1729) );
  AOI22X1TS U5495 ( .A0(mult2_out[9]), .A1(n4595), .B0(n4597), .B1(
        srmq_out[10]), .Y(n4577) );
  AOI22X1TS U5496 ( .A0(n1987), .A1(srmq_out[9]), .B0(n4592), .B1(srmq_out[8]), 
        .Y(n4576) );
  NAND2X1TS U5497 ( .A(n4577), .B(n4576), .Y(n1728) );
  AOI22X1TS U5498 ( .A0(n1987), .A1(srmq_out[8]), .B0(n4592), .B1(srmq_out[7]), 
        .Y(n4579) );
  AOI22X1TS U5499 ( .A0(mult2_out[8]), .A1(n4595), .B0(n4597), .B1(srmq_out[9]), .Y(n4578) );
  NAND2X1TS U5500 ( .A(n4579), .B(n4578), .Y(n1727) );
  AOI22X1TS U5501 ( .A0(n4592), .A1(srmq_out[6]), .B0(n4597), .B1(srmq_out[8]), 
        .Y(n4581) );
  AOI22X1TS U5502 ( .A0(mult2_out[7]), .A1(n4595), .B0(n1987), .B1(srmq_out[7]), .Y(n4580) );
  NAND2X1TS U5503 ( .A(n4581), .B(n4580), .Y(n1726) );
  AOI22X1TS U5504 ( .A0(mult2_out[6]), .A1(n4595), .B0(n4592), .B1(srmq_out[5]), .Y(n4583) );
  AOI22X1TS U5505 ( .A0(n1987), .A1(srmq_out[6]), .B0(n4597), .B1(srmq_out[7]), 
        .Y(n4582) );
  NAND2X1TS U5506 ( .A(n4583), .B(n4582), .Y(n1725) );
  AOI22X1TS U5507 ( .A0(mult2_out[5]), .A1(n4595), .B0(n1987), .B1(srmq_out[5]), .Y(n4585) );
  AOI22X1TS U5508 ( .A0(n4592), .A1(srmq_out[4]), .B0(n4597), .B1(srmq_out[6]), 
        .Y(n4584) );
  NAND2X1TS U5509 ( .A(n4585), .B(n4584), .Y(n1724) );
  AOI22X1TS U5510 ( .A0(n1987), .A1(srmq_out[4]), .B0(n4592), .B1(srmq_out[3]), 
        .Y(n4587) );
  AOI22X1TS U5511 ( .A0(mult2_out[4]), .A1(n4595), .B0(n4597), .B1(srmq_out[5]), .Y(n4586) );
  NAND2X1TS U5512 ( .A(n4587), .B(n4586), .Y(n1723) );
  AOI22X1TS U5513 ( .A0(mult2_out[3]), .A1(n4595), .B0(n1987), .B1(srmq_out[3]), .Y(n4589) );
  AOI22X1TS U5514 ( .A0(n4592), .A1(srmq_out[2]), .B0(n4597), .B1(srmq_out[4]), 
        .Y(n4588) );
  NAND2X1TS U5515 ( .A(n4589), .B(n4588), .Y(n1722) );
  AOI22X1TS U5516 ( .A0(mult2_out[2]), .A1(n4595), .B0(n4597), .B1(srmq_out[3]), .Y(n4591) );
  AOI22X1TS U5517 ( .A0(n1987), .A1(srmq_out[2]), .B0(n4592), .B1(srmq_out[1]), 
        .Y(n4590) );
  NAND2X1TS U5518 ( .A(n4591), .B(n4590), .Y(n1721) );
  AOI22X1TS U5519 ( .A0(n1987), .A1(srmq_out[1]), .B0(n4592), .B1(srmq_out[0]), 
        .Y(n4594) );
  AOI22X1TS U5520 ( .A0(mult2_out[1]), .A1(n4595), .B0(n4597), .B1(srmq_out[2]), .Y(n4593) );
  NAND2X1TS U5521 ( .A(n4594), .B(n4593), .Y(n1720) );
  AOI22X1TS U5522 ( .A0(n4595), .A1(mult2_out[0]), .B0(n1987), .B1(srmq_out[0]), .Y(n4596) );
  OAI2BB1X1TS U5523 ( .A0N(n4597), .A1N(srmq_out[1]), .B0(n4596), .Y(n1719) );
  AOI22X1TS U5524 ( .A0(n_input[31]), .A1(n4602), .B0(n4601), .B1(
        aluone_out[31]), .Y(n4600) );
  AOI22X1TS U5525 ( .A0(regres_out[31]), .A1(n4603), .B0(regres_out[30]), .B1(
        n4598), .Y(n4599) );
  NAND2X1TS U5526 ( .A(n4600), .B(n4599), .Y(n1718) );
  AOI22X1TS U5527 ( .A0(n4602), .A1(n_input[0]), .B0(n4601), .B1(aluone_out[0]), .Y(n4606) );
  AOI22X1TS U5528 ( .A0(regres_out[1]), .A1(n4604), .B0(regres_out[0]), .B1(
        n4603), .Y(n4605) );
  NAND2X1TS U5529 ( .A(n4606), .B(n4605), .Y(n1687) );
  OA21XLTS U5530 ( .A0(reg_i), .A1(regi_out[1]), .B0(n4607), .Y(n1685) );
  INVX2TS U5531 ( .A(reg_sp), .Y(n4609) );
  AOI22X1TS U5532 ( .A0(n4612), .A1(regsc_out), .B0(regsa_out), .B1(n4610), 
        .Y(n4608) );
  XNOR2X1TS U5533 ( .A(regsb_out), .B(n4608), .Y(n4611) );
  AO22XLTS U5534 ( .A0(n4609), .A1(regsp_out), .B0(reg_sp), .B1(n4611), .Y(
        n1683) );
  AO22XLTS U5535 ( .A0(n4612), .A1(n4611), .B0(n4610), .B1(regsq_out), .Y(
        n1682) );
  INVX2TS U5536 ( .A(reg_es0), .Y(n4632) );
  NOR3BX1TS U5537 ( .AN(mux7), .B(mux11), .C(n4632), .Y(n4627) );
  CLKAND2X2TS U5538 ( .A(mux11), .B(reg_es0), .Y(n4631) );
  AOI22X1TS U5539 ( .A0(reges_out[0]), .A1(n4627), .B0(n4631), .B1(
        aluone_out[0]), .Y(n4614) );
  NOR3X1TS U5540 ( .A(mux11), .B(mux7), .C(n4632), .Y(n4628) );
  AOI22X1TS U5541 ( .A0(reget_out[0]), .A1(n4628), .B0(reges0_out[0]), .B1(
        n4632), .Y(n4613) );
  NAND2X1TS U5542 ( .A(n4614), .B(n4613), .Y(n1681) );
  AOI22X1TS U5543 ( .A0(reget_out[1]), .A1(n4628), .B0(n4631), .B1(
        aluone_out[1]), .Y(n4616) );
  AOI22X1TS U5544 ( .A0(reges0_out[1]), .A1(n4632), .B0(reges_out[1]), .B1(
        n4627), .Y(n4615) );
  NAND2X1TS U5545 ( .A(n4616), .B(n4615), .Y(n1680) );
  AOI22X1TS U5546 ( .A0(reget_out[2]), .A1(n4628), .B0(n4631), .B1(
        aluone_out[2]), .Y(n4618) );
  AOI22X1TS U5547 ( .A0(reges_out[2]), .A1(n4627), .B0(reges0_out[2]), .B1(
        n4632), .Y(n4617) );
  NAND2X1TS U5548 ( .A(n4618), .B(n4617), .Y(n1679) );
  AOI22X1TS U5549 ( .A0(reget_out[3]), .A1(n4628), .B0(n4631), .B1(
        aluone_out[3]), .Y(n4620) );
  AOI22X1TS U5550 ( .A0(reges0_out[3]), .A1(n4632), .B0(reges_out[3]), .B1(
        n4627), .Y(n4619) );
  NAND2X1TS U5551 ( .A(n4620), .B(n4619), .Y(n1678) );
  AOI22X1TS U5552 ( .A0(reget_out[4]), .A1(n4628), .B0(n4631), .B1(
        aluone_out[4]), .Y(n4622) );
  AOI22X1TS U5553 ( .A0(reges_out[4]), .A1(n4627), .B0(reges0_out[4]), .B1(
        n4632), .Y(n4621) );
  NAND2X1TS U5554 ( .A(n4622), .B(n4621), .Y(n1677) );
  AOI22X1TS U5555 ( .A0(reget_out[5]), .A1(n4628), .B0(n4631), .B1(
        aluone_out[5]), .Y(n4624) );
  AOI22X1TS U5556 ( .A0(reges0_out[5]), .A1(n4632), .B0(reges_out[5]), .B1(
        n4627), .Y(n4623) );
  NAND2X1TS U5557 ( .A(n4624), .B(n4623), .Y(n1676) );
  AOI22X1TS U5558 ( .A0(reget_out[6]), .A1(n4628), .B0(n4631), .B1(
        aluone_out[6]), .Y(n4626) );
  AOI22X1TS U5559 ( .A0(reges_out[6]), .A1(n4627), .B0(reges0_out[6]), .B1(
        n4632), .Y(n4625) );
  NAND2X1TS U5560 ( .A(n4626), .B(n4625), .Y(n1675) );
  AOI22X1TS U5561 ( .A0(reges_out[7]), .A1(n4627), .B0(n4631), .B1(
        aluone_out[7]), .Y(n4630) );
  AOI22X1TS U5562 ( .A0(reges0_out[7]), .A1(n4632), .B0(reget_out[7]), .B1(
        n4628), .Y(n4629) );
  NAND2X1TS U5563 ( .A(n4630), .B(n4629), .Y(n1674) );
  AO22XLTS U5564 ( .A0(reges0_out[8]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[8]), .Y(n1673) );
  AO22XLTS U5565 ( .A0(reges0_out[9]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[9]), .Y(n1672) );
  AO22XLTS U5566 ( .A0(reges0_out[10]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[10]), .Y(n1671) );
  AO22XLTS U5567 ( .A0(reges0_out[11]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[11]), .Y(n1670) );
  AO22XLTS U5568 ( .A0(reges0_out[12]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[12]), .Y(n1669) );
  AO22XLTS U5569 ( .A0(reges0_out[13]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[13]), .Y(n1668) );
  AO22XLTS U5570 ( .A0(reges0_out[14]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[14]), .Y(n1667) );
  AO22XLTS U5571 ( .A0(reges0_out[15]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[15]), .Y(n1666) );
  AO22XLTS U5572 ( .A0(reges0_out[16]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[16]), .Y(n1665) );
  AO22XLTS U5573 ( .A0(reges0_out[17]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[17]), .Y(n1664) );
  AO22XLTS U5574 ( .A0(reges0_out[18]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[18]), .Y(n1663) );
  AO22XLTS U5575 ( .A0(reges0_out[19]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[19]), .Y(n1662) );
  AO22XLTS U5576 ( .A0(reges0_out[20]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[20]), .Y(n1661) );
  AO22XLTS U5577 ( .A0(reges0_out[21]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[21]), .Y(n1660) );
  AO22XLTS U5578 ( .A0(reges0_out[22]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[22]), .Y(n1659) );
  AO22XLTS U5579 ( .A0(reges0_out[23]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[23]), .Y(n1658) );
  AO22XLTS U5580 ( .A0(reges0_out[24]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[24]), .Y(n1657) );
  AO22XLTS U5581 ( .A0(reges0_out[25]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[25]), .Y(n1656) );
  AO22XLTS U5582 ( .A0(reges0_out[26]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[26]), .Y(n1655) );
  AO22XLTS U5583 ( .A0(reges0_out[27]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[27]), .Y(n1654) );
  AO22XLTS U5584 ( .A0(reges0_out[28]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[28]), .Y(n1653) );
  AO22XLTS U5585 ( .A0(reges0_out[29]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[29]), .Y(n1652) );
  AO22XLTS U5586 ( .A0(reges0_out[30]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[30]), .Y(n1651) );
  AO22XLTS U5588 ( .A0(reges0_out[31]), .A1(n4632), .B0(n4631), .B1(
        aluone_out[31]), .Y(n1649) );
  AOI211XLTS U5589 ( .A0(regres_out[5]), .A1(n4774), .B0(regres_out[31]), .C0(
        regres_out[30]), .Y(n4650) );
  NOR4XLTS U5590 ( .A(regres_out[29]), .B(regres_out[28]), .C(regres_out[27]), 
        .D(regres_out[26]), .Y(n4649) );
  NOR4XLTS U5591 ( .A(regres_out[9]), .B(regres_out[8]), .C(regres_out[7]), 
        .D(regres_out[6]), .Y(n4648) );
  NOR4XLTS U5592 ( .A(regres_out[21]), .B(regres_out[20]), .C(regres_out[19]), 
        .D(regres_out[18]), .Y(n4636) );
  NOR4XLTS U5593 ( .A(regres_out[25]), .B(regres_out[24]), .C(regres_out[23]), 
        .D(regres_out[22]), .Y(n4635) );
  NOR4XLTS U5594 ( .A(regres_out[13]), .B(regres_out[12]), .C(regres_out[11]), 
        .D(regres_out[10]), .Y(n4634) );
  NOR4XLTS U5595 ( .A(regres_out[17]), .B(regres_out[16]), .C(regres_out[15]), 
        .D(regres_out[14]), .Y(n4633) );
  NAND4XLTS U5596 ( .A(n4636), .B(n4635), .C(n4634), .D(n4633), .Y(n4646) );
  INVX2TS U5597 ( .A(regres_out[1]), .Y(n4638) );
  INVX2TS U5598 ( .A(regres_out[0]), .Y(n4637) );
  AOI211XLTS U5599 ( .A0(regindex_out[1]), .A1(n4638), .B0(regindex_out[0]), 
        .C0(n4637), .Y(n4640) );
  OAI22X1TS U5600 ( .A0(regindex_out[1]), .A1(n4638), .B0(regindex_out[2]), 
        .B1(n4642), .Y(n4639) );
  OAI22X1TS U5601 ( .A0(n4640), .A1(n4639), .B0(regres_out[3]), .B1(n4773), 
        .Y(n4641) );
  AOI21X1TS U5602 ( .A0(regindex_out[2]), .A1(n4642), .B0(n4641), .Y(n4645) );
  AO22XLTS U5603 ( .A0(n4784), .A1(regres_out[4]), .B0(n4773), .B1(
        regres_out[3]), .Y(n4644) );
  OA22X1TS U5604 ( .A0(n4784), .A1(regres_out[4]), .B0(n4774), .B1(
        regres_out[5]), .Y(n4643) );
  OAI32X1TS U5605 ( .A0(n4646), .A1(n4645), .A2(n4644), .B0(n4643), .B1(n4646), 
        .Y(n4647) );
  NAND4XLTS U5606 ( .A(n4650), .B(n4649), .C(n4648), .D(n4647), .Y(\comp2/N0 )
         );
  AOI22X1TS U5607 ( .A0(regcurrterm_out[24]), .A1(n4775), .B0(
        regcurrterm_out[25]), .B1(n4781), .Y(n4652) );
  OAI22X1TS U5608 ( .A0(regcurrterm_out[24]), .A1(n4775), .B0(
        regcurrterm_out[23]), .B1(n4785), .Y(n4651) );
  AOI22X1TS U5609 ( .A0(regsum_out[25]), .A1(n4787), .B0(n4652), .B1(n4651), 
        .Y(n4653) );
  AOI222XLTS U5610 ( .A0(regcurrterm_out[26]), .A1(n4653), .B0(
        regcurrterm_out[26]), .B1(n4782), .C0(n4653), .C1(n4782), .Y(n4654) );
  AOI222XLTS U5611 ( .A0(n4654), .A1(regsum_out[27]), .B0(n4654), .B1(n4808), 
        .C0(regsum_out[27]), .C1(n4808), .Y(n4655) );
  AOI21X1TS U5612 ( .A0(regcurrterm_out[28]), .A1(n4776), .B0(n4655), .Y(n4657) );
  OAI22X1TS U5613 ( .A0(regcurrterm_out[28]), .A1(n4776), .B0(
        regcurrterm_out[29]), .B1(n4786), .Y(n4656) );
  OAI22X1TS U5614 ( .A0(n4657), .A1(n4656), .B0(regsum_out[29]), .B1(n4805), 
        .Y(n4658) );
  AOI222XLTS U5615 ( .A0(regcurrterm_out[30]), .A1(n4783), .B0(
        regcurrterm_out[30]), .B1(n4658), .C0(n4783), .C1(n4658), .Y(
        \comp1/N0 ) );
  AOI32X1TS U5616 ( .A0(n4664), .A1(n4663), .A2(n4714), .B0(n4662), .B1(
        m17_out[30]), .Y(n4665) );
  AOI21X1TS U5617 ( .A0(n4667), .A1(n4666), .B0(n4665), .Y(n4668) );
  NAND2X1TS U5618 ( .A(n4669), .B(n4668), .Y(alutwo_out[30]) );
  AOI21X1TS U5619 ( .A0(n4672), .A1(n4671), .B0(n4670), .Y(n4682) );
  INVX2TS U5620 ( .A(n4673), .Y(n4675) );
  NAND2X1TS U5621 ( .A(n4679), .B(n4714), .Y(n4674) );
  OAI22X1TS U5622 ( .A0(n4682), .A1(n2456), .B0(n4681), .B1(n4680), .Y(
        alutwo_out[24]) );
  AOI22X1TS U5623 ( .A0(n4689), .A1(n4686), .B0(n4710), .B1(m17_out[16]), .Y(
        n4692) );
  AOI32X1TS U5624 ( .A0(n4693), .A1(m17_out[17]), .A2(n4692), .B0(n4691), .B1(
        n4690), .Y(n4694) );
  OA21XLTS U5625 ( .A0(n4699), .A1(n4698), .B0(n4697), .Y(n4707) );
  OAI22X1TS U5626 ( .A0(n4707), .A1(n2456), .B0(n4706), .B1(n4705), .Y(
        alutwo_out[13]) );
  OAI32X1TS U5627 ( .A0(n2456), .A1(n4713), .A2(n4712), .B0(n4711), .B1(n2456), 
        .Y(n4720) );
  OAI31X1TS U5628 ( .A0(n4717), .A1(n4716), .A2(n4715), .B0(n4714), .Y(n4719)
         );
  OAI32X1TS U5629 ( .A0(n4720), .A1(n4719), .A2(n4718), .B0(n4721), .B1(n4720), 
        .Y(n4723) );
  AOI32X1TS U5630 ( .A0(n4724), .A1(n4723), .A2(n4722), .B0(n4721), .B1(n4723), 
        .Y(alutwo_out[9]) );
  AOI22X1TS U5631 ( .A0(regcurrterm_out[27]), .A1(n4733), .B0(n4729), .B1(
        regacc_out[27]), .Y(n4728) );
  AOI22X1TS U5632 ( .A0(rf_aout[27]), .A1(n4732), .B0(n4731), .B1(
        regreg_out[27]), .Y(n4727) );
  OAI21XLTS U5633 ( .A0(reges0_out[4]), .A1(n4725), .B0(n4730), .Y(n4726) );
  NAND3XLTS U5634 ( .A(n4728), .B(n4727), .C(n4726), .Y(m2_out[27]) );
  AOI22X1TS U5635 ( .A0(reges0_out[1]), .A1(n4730), .B0(n4729), .B1(
        regacc_out[24]), .Y(n4736) );
  AOI22X1TS U5636 ( .A0(rf_aout[24]), .A1(n4732), .B0(n4731), .B1(
        regreg_out[24]), .Y(n4735) );
  OAI21XLTS U5637 ( .A0(regcurrterm_out[24]), .A1(mux2[0]), .B0(n4733), .Y(
        n4734) );
  NAND3XLTS U5638 ( .A(n4736), .B(n4735), .C(n4734), .Y(m2_out[24]) );
  AOI22X1TS U5639 ( .A0(n4740), .A1(alutwo_out[6]), .B0(n4739), .B1(
        regsum_out[29]), .Y(n4738) );
  AOI32X1TS U5640 ( .A0(n4743), .A1(n4738), .A2(n4737), .B0(n4741), .B1(n4738), 
        .Y(m3_out[29]) );
  AOI22X1TS U5641 ( .A0(n4740), .A1(alutwo_out[4]), .B0(n4739), .B1(
        regsum_out[27]), .Y(n4742) );
  INVX2TS U5642 ( .A(rf_aout[27]), .Y(n4748) );
  AOI32X1TS U5643 ( .A0(n4743), .A1(n4742), .A2(n4748), .B0(n4741), .B1(n4742), 
        .Y(m3_out[27]) );
  OAI21XLTS U5644 ( .A0(regsq_out), .A1(mux23), .B0(n3286), .Y(n4745) );
  AOI22X1TS U5645 ( .A0(n4771), .A1(rf_aout[31]), .B0(n4769), .B1(
        calculator_input[31]), .Y(n4744) );
  NAND2X1TS U5646 ( .A(n4745), .B(n4744), .Y(m14_out[31]) );
  OAI22X1TS U5647 ( .A0(n1991), .A1(alutwo_out[4]), .B0(calculator_input[27]), 
        .B1(n4746), .Y(n4747) );
  AOI22X1TS U5648 ( .A0(n4771), .A1(n4748), .B0(n4747), .B1(n4750), .Y(
        m14_out[27]) );
  INVX2TS U5649 ( .A(alutwo_out[1]), .Y(n4752) );
  OAI22X1TS U5650 ( .A0(rf_aout[24]), .A1(n4750), .B0(calculator_input[24]), 
        .B1(n4749), .Y(n4751) );
  AOI21X1TS U5651 ( .A0(n3286), .A1(n4752), .B0(n4751), .Y(m14_out[24]) );
  AOI22X1TS U5652 ( .A0(n3286), .A1(srmq_out[45]), .B0(n4769), .B1(
        calculator_input[22]), .Y(n4753) );
  OAI2BB1X1TS U5653 ( .A0N(n4771), .A1N(rf_aout[22]), .B0(n4753), .Y(
        m14_out[22]) );
  AOI22X1TS U5654 ( .A0(n3286), .A1(srmq_out[44]), .B0(n4769), .B1(
        calculator_input[21]), .Y(n4754) );
  OAI2BB1X1TS U5655 ( .A0N(n4771), .A1N(rf_aout[21]), .B0(n4754), .Y(
        m14_out[21]) );
  AOI22X1TS U5656 ( .A0(n3286), .A1(srmq_out[43]), .B0(n4769), .B1(
        calculator_input[20]), .Y(n4755) );
  OAI2BB1X1TS U5657 ( .A0N(n4771), .A1N(rf_aout[20]), .B0(n4755), .Y(
        m14_out[20]) );
  AOI22X1TS U5658 ( .A0(n3286), .A1(srmq_out[41]), .B0(n4769), .B1(
        calculator_input[18]), .Y(n4756) );
  OAI2BB1X1TS U5659 ( .A0N(n4771), .A1N(rf_aout[18]), .B0(n4756), .Y(
        m14_out[18]) );
  AOI22X1TS U5660 ( .A0(n3286), .A1(srmq_out[40]), .B0(n4769), .B1(
        calculator_input[17]), .Y(n4757) );
  OAI2BB1X1TS U5661 ( .A0N(n4771), .A1N(rf_aout[17]), .B0(n4757), .Y(
        m14_out[17]) );
  AOI22X1TS U5662 ( .A0(n3286), .A1(srmq_out[38]), .B0(n4769), .B1(
        calculator_input[15]), .Y(n4758) );
  OAI2BB1X1TS U5663 ( .A0N(n4771), .A1N(rf_aout[15]), .B0(n4758), .Y(
        m14_out[15]) );
  AOI22X1TS U5664 ( .A0(n3286), .A1(srmq_out[36]), .B0(n4769), .B1(
        calculator_input[13]), .Y(n4759) );
  OAI2BB1X1TS U5665 ( .A0N(n4771), .A1N(rf_aout[13]), .B0(n4759), .Y(
        m14_out[13]) );
  AOI22X1TS U5666 ( .A0(n3286), .A1(srmq_out[35]), .B0(n4769), .B1(
        calculator_input[12]), .Y(n4760) );
  OAI2BB1X1TS U5667 ( .A0N(n4771), .A1N(rf_aout[12]), .B0(n4760), .Y(
        m14_out[12]) );
  AOI22X1TS U5668 ( .A0(n3286), .A1(srmq_out[34]), .B0(n4769), .B1(
        calculator_input[11]), .Y(n4761) );
  OAI2BB1X1TS U5669 ( .A0N(n4771), .A1N(rf_aout[11]), .B0(n4761), .Y(
        m14_out[11]) );
  AOI22X1TS U5670 ( .A0(n3286), .A1(srmq_out[33]), .B0(n4769), .B1(
        calculator_input[10]), .Y(n4762) );
  OAI2BB1X1TS U5671 ( .A0N(n4771), .A1N(rf_aout[10]), .B0(n4762), .Y(
        m14_out[10]) );
  AOI22X1TS U5672 ( .A0(n3286), .A1(srmq_out[30]), .B0(n4769), .B1(
        calculator_input[7]), .Y(n4763) );
  OAI2BB1X1TS U5673 ( .A0N(n4771), .A1N(rf_aout[7]), .B0(n4763), .Y(m14_out[7]) );
  AOI22X1TS U5674 ( .A0(n3286), .A1(srmq_out[29]), .B0(n4769), .B1(
        calculator_input[6]), .Y(n4764) );
  OAI2BB1X1TS U5675 ( .A0N(n4771), .A1N(rf_aout[6]), .B0(n4764), .Y(m14_out[6]) );
  AOI22X1TS U5676 ( .A0(n3286), .A1(srmq_out[28]), .B0(n4769), .B1(
        calculator_input[5]), .Y(n4765) );
  OAI2BB1X1TS U5677 ( .A0N(n4771), .A1N(rf_aout[5]), .B0(n4765), .Y(m14_out[5]) );
  AOI22X1TS U5678 ( .A0(n3286), .A1(srmq_out[26]), .B0(n4769), .B1(
        calculator_input[3]), .Y(n4766) );
  OAI2BB1X1TS U5679 ( .A0N(n4771), .A1N(rf_aout[3]), .B0(n4766), .Y(m14_out[3]) );
  AOI22X1TS U5680 ( .A0(n3286), .A1(srmq_out[25]), .B0(n4769), .B1(
        calculator_input[2]), .Y(n4767) );
  OAI2BB1X1TS U5681 ( .A0N(n4771), .A1N(rf_aout[2]), .B0(n4767), .Y(m14_out[2]) );
  AOI22X1TS U5682 ( .A0(n3286), .A1(srmq_out[24]), .B0(n4769), .B1(
        calculator_input[1]), .Y(n4768) );
  OAI2BB1X1TS U5683 ( .A0N(n4771), .A1N(rf_aout[1]), .B0(n4768), .Y(m14_out[1]) );
  AOI22X1TS U5684 ( .A0(n3286), .A1(srmq_out[23]), .B0(n4769), .B1(
        calculator_input[0]), .Y(n4770) );
  OAI2BB1X1TS U5685 ( .A0N(n4771), .A1N(rf_aout[0]), .B0(n4770), .Y(m14_out[0]) );
endmodule

